//
// Copyright (C) 2014, 2017-2018 Chris McClelland
//
// Permission is hereby granted, free of charge, to any person obtaining a copy of this software
// and associated documentation files (the "Software"), to deal in the Software without
// restriction, including without limitation the rights to use, copy, modify, merge, publish,
// distribute, sublicense, and/or sell copies of the Software, and to permit persons to whom the
// Software is furnished to do so, subject to the following conditions:
//
// The above copyright  notice and this permission notice  shall be included in all copies or
// substantial portions of the Software.
//
// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR IMPLIED, INCLUDING
// BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND
// NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM,
// DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE SOFTWARE.
//
module pcie_sv(
    // Clock, resets, PCIe physical RX & TX
    input logic pcieRefClk_in,
    input logic pcieNPOR_in,
    input logic pciePERST_in,
    input logic[3:0] pcieRX_in,
    output logic[3:0] pcieTX_out,

    // Application interface
    output logic pcieClk_out,
    output tlp_xcvr_pkg::BusID cfgBusDev_out,

    output tlp_xcvr_pkg::uint64 rxData_out,
    output logic rxSOP_out,
    output logic rxEOP_out,
    output logic rxValid_out,
    input logic rxReady_in,

    input tlp_xcvr_pkg::uint64 txData_in,
    input logic txSOP_in,
    input logic txEOP_in,
    input logic txValid_in,
    output logic txReady_out,

    // Control & Pipe signals for simulation connection
    input  wire [31:0] hip_ctrl_test_in,          //   hip_ctrl.test_in
    input  wire        hip_ctrl_simu_mode_pipe,   //           .simu_mode_pipe
    input  wire        hip_pipe_sim_pipe_pclk_in, //   hip_pipe.sim_pipe_pclk_in
    output wire [1:0]  hip_pipe_sim_pipe_rate,    //           .sim_pipe_rate
    output wire [4:0]  hip_pipe_sim_ltssmstate,   //           .sim_ltssmstate
    output wire [2:0]  hip_pipe_eidleinfersel0,   //           .eidleinfersel0
    output wire [2:0]  hip_pipe_eidleinfersel1,   //           .eidleinfersel1
    output wire [2:0]  hip_pipe_eidleinfersel2,   //           .eidleinfersel2
    output wire [2:0]  hip_pipe_eidleinfersel3,   //           .eidleinfersel3
    output wire [1:0]  hip_pipe_powerdown0,       //           .powerdown0
    output wire [1:0]  hip_pipe_powerdown1,       //           .powerdown1
    output wire [1:0]  hip_pipe_powerdown2,       //           .powerdown2
    output wire [1:0]  hip_pipe_powerdown3,       //           .powerdown3
    output wire        hip_pipe_rxpolarity0,      //           .rxpolarity0
    output wire        hip_pipe_rxpolarity1,      //           .rxpolarity1
    output wire        hip_pipe_rxpolarity2,      //           .rxpolarity2
    output wire        hip_pipe_rxpolarity3,      //           .rxpolarity3
    output wire        hip_pipe_txcompl0,         //           .txcompl0
    output wire        hip_pipe_txcompl1,         //           .txcompl1
    output wire        hip_pipe_txcompl2,         //           .txcompl2
    output wire        hip_pipe_txcompl3,         //           .txcompl3
    output wire [7:0]  hip_pipe_txdata0,          //           .txdata0
    output wire [7:0]  hip_pipe_txdata1,          //           .txdata1
    output wire [7:0]  hip_pipe_txdata2,          //           .txdata2
    output wire [7:0]  hip_pipe_txdata3,          //           .txdata3
    output wire        hip_pipe_txdatak0,         //           .txdatak0
    output wire        hip_pipe_txdatak1,         //           .txdatak1
    output wire        hip_pipe_txdatak2,         //           .txdatak2
    output wire        hip_pipe_txdatak3,         //           .txdatak3
    output wire        hip_pipe_txdetectrx0,      //           .txdetectrx0
    output wire        hip_pipe_txdetectrx1,      //           .txdetectrx1
    output wire        hip_pipe_txdetectrx2,      //           .txdetectrx2
    output wire        hip_pipe_txdetectrx3,      //           .txdetectrx3
    output wire        hip_pipe_txelecidle0,      //           .txelecidle0
    output wire        hip_pipe_txelecidle1,      //           .txelecidle1
    output wire        hip_pipe_txelecidle2,      //           .txelecidle2
    output wire        hip_pipe_txelecidle3,      //           .txelecidle3
    output wire        hip_pipe_txdeemph0,        //           .txdeemph0
    output wire        hip_pipe_txdeemph1,        //           .txdeemph1
    output wire        hip_pipe_txdeemph2,        //           .txdeemph2
    output wire        hip_pipe_txdeemph3,        //           .txdeemph3
    output wire [2:0]  hip_pipe_txmargin0,        //           .txmargin0
    output wire [2:0]  hip_pipe_txmargin1,        //           .txmargin1
    output wire [2:0]  hip_pipe_txmargin2,        //           .txmargin2
    output wire [2:0]  hip_pipe_txmargin3,        //           .txmargin3
    output wire        hip_pipe_txswing0,         //           .txswing0
    output wire        hip_pipe_txswing1,         //           .txswing1
    output wire        hip_pipe_txswing2,         //           .txswing2
    output wire        hip_pipe_txswing3,         //           .txswing3
    input  wire        hip_pipe_phystatus0,       //           .phystatus0
    input  wire        hip_pipe_phystatus1,       //           .phystatus1
    input  wire        hip_pipe_phystatus2,       //           .phystatus2
    input  wire        hip_pipe_phystatus3,       //           .phystatus3
    input  wire [7:0]  hip_pipe_rxdata0,          //           .rxdata0
    input  wire [7:0]  hip_pipe_rxdata1,          //           .rxdata1
    input  wire [7:0]  hip_pipe_rxdata2,          //           .rxdata2
    input  wire [7:0]  hip_pipe_rxdata3,          //           .rxdata3
    input  wire        hip_pipe_rxdatak0,         //           .rxdatak0
    input  wire        hip_pipe_rxdatak1,         //           .rxdatak1
    input  wire        hip_pipe_rxdatak2,         //           .rxdatak2
    input  wire        hip_pipe_rxdatak3,         //           .rxdatak3
    input  wire        hip_pipe_rxelecidle0,      //           .rxelecidle0
    input  wire        hip_pipe_rxelecidle1,      //           .rxelecidle1
    input  wire        hip_pipe_rxelecidle2,      //           .rxelecidle2
    input  wire        hip_pipe_rxelecidle3,      //           .rxelecidle3
    input  wire [2:0]  hip_pipe_rxstatus0,        //           .rxstatus0
    input  wire [2:0]  hip_pipe_rxstatus1,        //           .rxstatus1
    input  wire [2:0]  hip_pipe_rxstatus2,        //           .rxstatus2
    input  wire [2:0]  hip_pipe_rxstatus3,        //           .rxstatus3
    input  wire        hip_pipe_rxvalid0,         //           .rxvalid0
    input  wire        hip_pipe_rxvalid1,         //           .rxvalid1
    input  wire        hip_pipe_rxvalid2,         //           .rxvalid2
    input  wire        hip_pipe_rxvalid3          //           .rxvalid3
  );

  // Interconnect signals
  logic       pcieClk;
  logic       pllLocked;
  logic[3:0]  tl_cfg_add;
  logic[31:0] tl_cfg_ctl;
  logic[65:0] fiData;
  logic       fiValid;
  logic[65:0] foData;
  logic       foValid;
  logic       foReady;

  // Instantiate the Verilog config-region sampler unit provided by Altera
  altpcierd_tl_cfg_sample sampler(
    .pld_clk        (pcieClk),
    .rstn           (1'b1),
    .tl_cfg_add     (tl_cfg_add),
    .tl_cfg_ctl     (tl_cfg_ctl),
    .tl_cfg_ctl_wr  (1'b0),
    .tl_cfg_sts     ('0),
    .tl_cfg_sts_wr  (1'b0),
    .cfg_busdev     (cfgBusDev_out[15:3])  // 13-bit device ID assigned to the FPGA on enumeration
  );
  assign cfgBusDev_out[2:0] = 0;

  // Small FIFO to avoid rxData being lost because of the two-clock latency from the PCIe IP.
  buffer_fifo#(
    .WIDTH           (66),    // space for 64-bit data word and the SOP & EOP flags
    .DEPTH           (2),     // space for four entries
    .BLOCK_RAM       (0)      // just use regular registers
  ) recv_fifo (
    .clk_in          (pcieClk),
    .reset_in        (),
    .depth_out       (),

    // Producer end
    .iData_in        (fiData),
    .iValid_in       (fiValid),
    .iReady_out      (),
    .iReadyChunk_out (),

    // Consumer end
    .oData_out       (foData),
    .oValid_out      (foValid),
    .oReady_in       (foReady),
    .oValidChunk_out ()
  );

  // Drive pcieClk externally
  assign pcieClk_out = pcieClk;

  // External connection to FIFO output
  assign rxData_out = foData[63:0];
  assign rxSOP_out = foData[64];
  assign rxEOP_out = foData[65];
  assign rxValid_out = foValid;
  assign foReady = rxReady_in;

  // The actual PCIe IP block
  altpcie_sv_hip_ast_hwtcl #(
    .ACDS_VERSION_HWTCL                       ("16.1"),
    .lane_mask_hwtcl                          ("x4"),
    .gen123_lane_rate_mode_hwtcl              ("Gen1 (2.5 Gbps)"),
    .port_type_hwtcl                          ("Native endpoint"),
    .pcie_spec_version_hwtcl                  ("2.1"),
    .ast_width_hwtcl                          ("Avalon-ST 64-bit"),
    .pll_refclk_freq_hwtcl                    ("100 MHz"),
    .set_pld_clk_x1_625MHz_hwtcl              (0),
    .use_ast_parity                           (0),
    .multiple_packets_per_cycle_hwtcl         (0),
    .in_cvp_mode_hwtcl                        (0),
    .use_pci_ext_hwtcl                        (0),
    .use_pcie_ext_hwtcl                       (0),
    .use_config_bypass_hwtcl                  (0),
    .enable_tl_only_sim_hwtcl                 (0),
    .hip_reconfig_hwtcl                       (0),
    .hip_tag_checking_hwtcl                   (1),
    .enable_power_on_rst_pulse_hwtcl          (0),
    .enable_pcisigtest_hwtcl                  (0),
    .bar0_size_mask_hwtcl                     (tlp_xcvr_pkg::BAR0_OFFSET_NBITS),
    .bar0_io_space_hwtcl                      ("Disabled"),
    .bar0_64bit_mem_space_hwtcl               ("Disabled"),
    .bar0_prefetchable_hwtcl                  ("Disabled"),
    .bar1_size_mask_hwtcl                     (0),
    .bar1_io_space_hwtcl                      ("Disabled"),
    .bar1_prefetchable_hwtcl                  ("Disabled"),
    .bar2_size_mask_hwtcl                     (tlp_xcvr_pkg::BAR0_OFFSET_NBITS),
    .bar2_io_space_hwtcl                      ("Disabled"),
    .bar2_64bit_mem_space_hwtcl               ("Enabled"),
    .bar2_prefetchable_hwtcl                  ("Enabled"),
    .bar3_size_mask_hwtcl                     (0),
    .bar3_io_space_hwtcl                      ("Disabled"),
    .bar3_prefetchable_hwtcl                  ("Disabled"),
    .bar4_size_mask_hwtcl                     (0),
    .bar4_io_space_hwtcl                      ("Disabled"),
    .bar4_64bit_mem_space_hwtcl               ("Disabled"),
    .bar4_prefetchable_hwtcl                  ("Disabled"),
    .bar5_size_mask_hwtcl                     (0),
    .bar5_io_space_hwtcl                      ("Disabled"),
    .bar5_prefetchable_hwtcl                  ("Disabled"),
    .expansion_base_address_register_hwtcl    (0),
    .io_window_addr_width_hwtcl               (0),
    .prefetchable_mem_window_addr_width_hwtcl (0),
    .vendor_id_hwtcl                          (4466),
    .device_id_hwtcl                          (57345),
    .revision_id_hwtcl                        (1),
    .class_code_hwtcl                         (16711680),
    .subsystem_vendor_id_hwtcl                (4466),
    .subsystem_device_id_hwtcl                (57345),
    .max_payload_size_hwtcl                   (256),
    .extend_tag_field_hwtcl                   ("32"),
    .completion_timeout_hwtcl                 ("ABCD"),
    .enable_completion_timeout_disable_hwtcl  (1),
    .use_aer_hwtcl                            (0),
    .ecrc_check_capable_hwtcl                 (0),
    .ecrc_gen_capable_hwtcl                   (0),
    .use_crc_forwarding_hwtcl                 (0),
    .port_link_number_hwtcl                   (1),
    .dll_active_report_support_hwtcl          (0),
    .surprise_down_error_support_hwtcl        (0),
    .slotclkcfg_hwtcl                         (1),
    .msi_multi_message_capable_hwtcl          ("4"),
    .msi_64bit_addressing_capable_hwtcl       ("true"),
    .msi_masking_capable_hwtcl                ("false"),
    .msi_support_hwtcl                        ("true"),
    .enable_function_msix_support_hwtcl       (0),
    .msix_table_size_hwtcl                    (0),
    .msix_table_offset_hwtcl                  ("0"),
    .msix_table_bir_hwtcl                     (0),
    .msix_pba_offset_hwtcl                    ("0"),
    .msix_pba_bir_hwtcl                       (0),
    .enable_slot_register_hwtcl               (0),
    .slot_power_scale_hwtcl                   (0),
    .slot_power_limit_hwtcl                   (0),
    .slot_number_hwtcl                        (0),
    .endpoint_l0_latency_hwtcl                (0),
    .endpoint_l1_latency_hwtcl                (0),
    .vsec_id_hwtcl                            (40960),
    .vsec_rev_hwtcl                           (0),
    .user_id_hwtcl                            (0),
    .millisecond_cycle_count_hwtcl            (124250),
    .port_width_be_hwtcl                      (8),
    .port_width_data_hwtcl                    (64),
    .gen3_dcbal_en_hwtcl                      (1),
    .enable_pipe32_sim_hwtcl                  (0),
    .fixed_preset_on                          (0),
    .bypass_cdc_hwtcl                         ("false"),
    .enable_rx_buffer_checking_hwtcl          ("false"),
    .disable_link_x2_support_hwtcl            ("false"),
    .wrong_device_id_hwtcl                    ("disable"),
    .data_pack_rx_hwtcl                       ("disable"),
    .ltssm_1ms_timeout_hwtcl                  ("disable"),
    .ltssm_freqlocked_check_hwtcl             ("disable"),
    .deskew_comma_hwtcl                       ("skp_eieos_deskw"),
    .device_number_hwtcl                      (0),
    .pipex1_debug_sel_hwtcl                   ("disable"),
    .pclk_out_sel_hwtcl                       ("pclk"),
    .no_soft_reset_hwtcl                      ("false"),
    .maximum_current_hwtcl                    (0),
    .d1_support_hwtcl                         ("false"),
    .d2_support_hwtcl                         ("false"),
    .d0_pme_hwtcl                             ("false"),
    .d1_pme_hwtcl                             ("false"),
    .d2_pme_hwtcl                             ("false"),
    .d3_hot_pme_hwtcl                         ("false"),
    .d3_cold_pme_hwtcl                        ("false"),
    .low_priority_vc_hwtcl                    ("single_vc"),
    .disable_snoop_packet_hwtcl               ("false"),
    .enable_l1_aspm_hwtcl                     ("false"),
    .rx_ei_l0s_hwtcl                          (0),
    .enable_l0s_aspm_hwtcl                    ("false"),
    .aspm_config_management_hwtcl             ("true"),
    .l1_exit_latency_sameclock_hwtcl          (0),
    .l1_exit_latency_diffclock_hwtcl          (0),
    .hot_plug_support_hwtcl                   (0),
    .extended_tag_reset_hwtcl                 ("false"),
    .no_command_completed_hwtcl               ("false"),
    .interrupt_pin_hwtcl                      ("inta"),
    .bridge_port_vga_enable_hwtcl             ("false"),
    .bridge_port_ssid_support_hwtcl           ("false"),
    .ssvid_hwtcl                              (0),
    .ssid_hwtcl                               (0),
    .eie_before_nfts_count_hwtcl              (4),
    .gen2_diffclock_nfts_count_hwtcl          (255),
    .gen2_sameclock_nfts_count_hwtcl          (255),
    .l0_exit_latency_sameclock_hwtcl          (6),
    .l0_exit_latency_diffclock_hwtcl          (6),
    .atomic_op_routing_hwtcl                  ("false"),
    .atomic_op_completer_32bit_hwtcl          ("false"),
    .atomic_op_completer_64bit_hwtcl          ("false"),
    .cas_completer_128bit_hwtcl               ("false"),
    .ltr_mechanism_hwtcl                      ("false"),
    .tph_completer_hwtcl                      ("false"),
    .extended_format_field_hwtcl              ("false"),
    .atomic_malformed_hwtcl                   ("true"),
    .flr_capability_hwtcl                     ("false"),
    .enable_adapter_half_rate_mode_hwtcl      ("false"),
    .vc0_clk_enable_hwtcl                     ("true"),
    .register_pipe_signals_hwtcl              ("false"),
    .skp_os_gen3_count_hwtcl                  (0),
    .tx_cdc_almost_empty_hwtcl                (5),
    .rx_l0s_count_idl_hwtcl                   (0),
    .cdc_dummy_insert_limit_hwtcl             (11),
    .ei_delay_powerdown_count_hwtcl           (10),
    .skp_os_schedule_count_hwtcl              (0),
    .fc_init_timer_hwtcl                      (1024),
    .l01_entry_latency_hwtcl                  (31),
    .flow_control_update_count_hwtcl          (30),
    .flow_control_timeout_count_hwtcl         (200),
    .retry_buffer_last_active_address_hwtcl   (2047),
    .reserved_debug_hwtcl                     (0),
    .bypass_clk_switch_hwtcl                  ("false"),
    .l2_async_logic_hwtcl                     ("disable"),
    .indicator_hwtcl                          (0),
    .diffclock_nfts_count_hwtcl               (128),
    .sameclock_nfts_count_hwtcl               (128),
    .rx_cdc_almost_full_hwtcl                 (12),
    .tx_cdc_almost_full_hwtcl                 (11),
    .credit_buffer_allocation_aux_hwtcl       ("absolute"),
    .vc0_rx_flow_ctrl_posted_header_hwtcl     (16),
    .vc0_rx_flow_ctrl_posted_data_hwtcl       (16),
    .vc0_rx_flow_ctrl_nonposted_header_hwtcl  (16),
    .vc0_rx_flow_ctrl_nonposted_data_hwtcl    (0),
    .vc0_rx_flow_ctrl_compl_header_hwtcl      (0),
    .vc0_rx_flow_ctrl_compl_data_hwtcl        (0),
    .cpl_spc_header_hwtcl                     (195),
    .cpl_spc_data_hwtcl                       (781),
    .gen3_rxfreqlock_counter_hwtcl            (0),
    .gen3_skip_ph2_ph3_hwtcl                  (0),
    .g3_bypass_equlz_hwtcl                    (0),
    .cvp_data_compressed_hwtcl                ("false"),
    .cvp_data_encrypted_hwtcl                 ("false"),
    .cvp_mode_reset_hwtcl                     ("false"),
    .cvp_clk_reset_hwtcl                      ("false"),
    .cseb_cpl_status_during_cvp_hwtcl         ("completer_abort"),
    .core_clk_sel_hwtcl                       ("core_clk_250"),
    .cvp_rate_sel_hwtcl                       ("full_rate"),
    .g3_dis_rx_use_prst_hwtcl                 ("true"),
    .g3_dis_rx_use_prst_ep_hwtcl              ("true"),
    .deemphasis_enable_hwtcl                  ("false"),
    .reconfig_to_xcvr_width                   (350),
    .reconfig_from_xcvr_width                 (230),
    .single_rx_detect_hwtcl                   (4),
    .hip_hard_reset_hwtcl                     (1),
    .use_cvp_update_core_pof_hwtcl            (0),
    .pcie_inspector_hwtcl                     (0),
    .tlp_inspector_hwtcl                      (1),
    .tlp_inspector_use_signal_probe_hwtcl     (0),
    .tlp_insp_trg_dw0_hwtcl                   (2049),
    .tlp_insp_trg_dw1_hwtcl                   (0),
    .tlp_insp_trg_dw2_hwtcl                   (0),
    .tlp_insp_trg_dw3_hwtcl                   (0),
    .hwtcl_override_g2_txvod                  (0),
    .rpre_emph_a_val_hwtcl                    (9),
    .rpre_emph_b_val_hwtcl                    (0),
    .rpre_emph_c_val_hwtcl                    (16),
    .rpre_emph_d_val_hwtcl                    (13),
    .rpre_emph_e_val_hwtcl                    (5),
    .rvod_sel_a_val_hwtcl                     (42),
    .rvod_sel_b_val_hwtcl                     (38),
    .rvod_sel_c_val_hwtcl                     (38),
    .rvod_sel_d_val_hwtcl                     (43),
    .rvod_sel_e_val_hwtcl                     (15),
    .hwtcl_override_g3rxcoef                  (0),
    .gen3_coeff_1_hwtcl                       (7),
    .gen3_coeff_1_sel_hwtcl                   ("preset_1"),
    .gen3_coeff_1_preset_hint_hwtcl           (0),
    .gen3_coeff_1_nxtber_more_ptr_hwtcl       (1),
    .gen3_coeff_1_nxtber_more_hwtcl           ("g3_coeff_1_nxtber_more"),
    .gen3_coeff_1_nxtber_less_ptr_hwtcl       (1),
    .gen3_coeff_1_nxtber_less_hwtcl           ("g3_coeff_1_nxtber_less"),
    .gen3_coeff_1_reqber_hwtcl                (0),
    .gen3_coeff_1_ber_meas_hwtcl              (2),
    .gen3_coeff_2_hwtcl                       (0),
    .gen3_coeff_2_sel_hwtcl                   ("preset_2"),
    .gen3_coeff_2_preset_hint_hwtcl           (0),
    .gen3_coeff_2_nxtber_more_ptr_hwtcl       (0),
    .gen3_coeff_2_nxtber_more_hwtcl           ("g3_coeff_2_nxtber_more"),
    .gen3_coeff_2_nxtber_less_ptr_hwtcl       (0),
    .gen3_coeff_2_nxtber_less_hwtcl           ("g3_coeff_2_nxtber_less"),
    .gen3_coeff_2_reqber_hwtcl                (0),
    .gen3_coeff_2_ber_meas_hwtcl              (0),
    .gen3_coeff_3_hwtcl                       (0),
    .gen3_coeff_3_sel_hwtcl                   ("preset_3"),
    .gen3_coeff_3_preset_hint_hwtcl           (0),
    .gen3_coeff_3_nxtber_more_ptr_hwtcl       (0),
    .gen3_coeff_3_nxtber_more_hwtcl           ("g3_coeff_3_nxtber_more"),
    .gen3_coeff_3_nxtber_less_ptr_hwtcl       (0),
    .gen3_coeff_3_nxtber_less_hwtcl           ("g3_coeff_3_nxtber_less"),
    .gen3_coeff_3_reqber_hwtcl                (0),
    .gen3_coeff_3_ber_meas_hwtcl              (0),
    .gen3_coeff_4_hwtcl                       (0),
    .gen3_coeff_4_sel_hwtcl                   ("preset_4"),
    .gen3_coeff_4_preset_hint_hwtcl           (0),
    .gen3_coeff_4_nxtber_more_ptr_hwtcl       (0),
    .gen3_coeff_4_nxtber_more_hwtcl           ("g3_coeff_4_nxtber_more"),
    .gen3_coeff_4_nxtber_less_ptr_hwtcl       (0),
    .gen3_coeff_4_nxtber_less_hwtcl           ("g3_coeff_4_nxtber_less"),
    .gen3_coeff_4_reqber_hwtcl                (0),
    .gen3_coeff_4_ber_meas_hwtcl              (0),
    .gen3_coeff_5_hwtcl                       (0),
    .gen3_coeff_5_sel_hwtcl                   ("preset_5"),
    .gen3_coeff_5_preset_hint_hwtcl           (0),
    .gen3_coeff_5_nxtber_more_ptr_hwtcl       (0),
    .gen3_coeff_5_nxtber_more_hwtcl           ("g3_coeff_5_nxtber_more"),
    .gen3_coeff_5_nxtber_less_ptr_hwtcl       (0),
    .gen3_coeff_5_nxtber_less_hwtcl           ("g3_coeff_5_nxtber_less"),
    .gen3_coeff_5_reqber_hwtcl                (0),
    .gen3_coeff_5_ber_meas_hwtcl              (0),
    .gen3_coeff_6_hwtcl                       (0),
    .gen3_coeff_6_sel_hwtcl                   ("preset_6"),
    .gen3_coeff_6_preset_hint_hwtcl           (0),
    .gen3_coeff_6_nxtber_more_ptr_hwtcl       (0),
    .gen3_coeff_6_nxtber_more_hwtcl           ("g3_coeff_6_nxtber_more"),
    .gen3_coeff_6_nxtber_less_ptr_hwtcl       (0),
    .gen3_coeff_6_nxtber_less_hwtcl           ("g3_coeff_6_nxtber_less"),
    .gen3_coeff_6_reqber_hwtcl                (0),
    .gen3_coeff_6_ber_meas_hwtcl              (0),
    .gen3_coeff_7_hwtcl                       (0),
    .gen3_coeff_7_sel_hwtcl                   ("preset_7"),
    .gen3_coeff_7_preset_hint_hwtcl           (0),
    .gen3_coeff_7_nxtber_more_ptr_hwtcl       (0),
    .gen3_coeff_7_nxtber_more_hwtcl           ("g3_coeff_7_nxtber_more"),
    .gen3_coeff_7_nxtber_less_ptr_hwtcl       (0),
    .gen3_coeff_7_nxtber_less_hwtcl           ("g3_coeff_7_nxtber_less"),
    .gen3_coeff_7_reqber_hwtcl                (0),
    .gen3_coeff_7_ber_meas_hwtcl              (0),
    .gen3_coeff_8_hwtcl                       (0),
    .gen3_coeff_8_sel_hwtcl                   ("preset_8"),
    .gen3_coeff_8_preset_hint_hwtcl           (0),
    .gen3_coeff_8_nxtber_more_ptr_hwtcl       (0),
    .gen3_coeff_8_nxtber_more_hwtcl           ("g3_coeff_8_nxtber_more"),
    .gen3_coeff_8_nxtber_less_ptr_hwtcl       (0),
    .gen3_coeff_8_nxtber_less_hwtcl           ("g3_coeff_8_nxtber_less"),
    .gen3_coeff_8_reqber_hwtcl                (0),
    .gen3_coeff_8_ber_meas_hwtcl              (0),
    .gen3_coeff_9_hwtcl                       (0),
    .gen3_coeff_9_sel_hwtcl                   ("preset_9"),
    .gen3_coeff_9_preset_hint_hwtcl           (0),
    .gen3_coeff_9_nxtber_more_ptr_hwtcl       (0),
    .gen3_coeff_9_nxtber_more_hwtcl           ("g3_coeff_9_nxtber_more"),
    .gen3_coeff_9_nxtber_less_ptr_hwtcl       (0),
    .gen3_coeff_9_nxtber_less_hwtcl           ("g3_coeff_9_nxtber_less"),
    .gen3_coeff_9_reqber_hwtcl                (0),
    .gen3_coeff_9_ber_meas_hwtcl              (0),
    .gen3_coeff_10_hwtcl                      (0),
    .gen3_coeff_10_sel_hwtcl                  ("preset_10"),
    .gen3_coeff_10_preset_hint_hwtcl          (0),
    .gen3_coeff_10_nxtber_more_ptr_hwtcl      (0),
    .gen3_coeff_10_nxtber_more_hwtcl          ("g3_coeff_10_nxtber_more"),
    .gen3_coeff_10_nxtber_less_ptr_hwtcl      (0),
    .gen3_coeff_10_nxtber_less_hwtcl          ("g3_coeff_10_nxtber_less"),
    .gen3_coeff_10_reqber_hwtcl               (0),
    .gen3_coeff_10_ber_meas_hwtcl             (0),
    .gen3_coeff_11_hwtcl                      (0),
    .gen3_coeff_11_sel_hwtcl                  ("preset_11"),
    .gen3_coeff_11_preset_hint_hwtcl          (0),
    .gen3_coeff_11_nxtber_more_ptr_hwtcl      (0),
    .gen3_coeff_11_nxtber_more_hwtcl          ("g3_coeff_11_nxtber_more"),
    .gen3_coeff_11_nxtber_less_ptr_hwtcl      (0),
    .gen3_coeff_11_nxtber_less_hwtcl          ("g3_coeff_11_nxtber_less"),
    .gen3_coeff_11_reqber_hwtcl               (0),
    .gen3_coeff_11_ber_meas_hwtcl             (0),
    .gen3_coeff_12_hwtcl                      (0),
    .gen3_coeff_12_sel_hwtcl                  ("preset_12"),
    .gen3_coeff_12_preset_hint_hwtcl          (0),
    .gen3_coeff_12_nxtber_more_ptr_hwtcl      (0),
    .gen3_coeff_12_nxtber_more_hwtcl          ("g3_coeff_12_nxtber_more"),
    .gen3_coeff_12_nxtber_less_ptr_hwtcl      (0),
    .gen3_coeff_12_nxtber_less_hwtcl          ("g3_coeff_12_nxtber_less"),
    .gen3_coeff_12_reqber_hwtcl               (0),
    .gen3_coeff_12_ber_meas_hwtcl             (0),
    .gen3_coeff_13_hwtcl                      (0),
    .gen3_coeff_13_sel_hwtcl                  ("preset_13"),
    .gen3_coeff_13_preset_hint_hwtcl          (0),
    .gen3_coeff_13_nxtber_more_ptr_hwtcl      (0),
    .gen3_coeff_13_nxtber_more_hwtcl          ("g3_coeff_13_nxtber_more"),
    .gen3_coeff_13_nxtber_less_ptr_hwtcl      (0),
    .gen3_coeff_13_nxtber_less_hwtcl          ("g3_coeff_13_nxtber_less"),
    .gen3_coeff_13_reqber_hwtcl               (0),
    .gen3_coeff_13_ber_meas_hwtcl             (0),
    .gen3_coeff_14_hwtcl                      (0),
    .gen3_coeff_14_sel_hwtcl                  ("preset_14"),
    .gen3_coeff_14_preset_hint_hwtcl          (0),
    .gen3_coeff_14_nxtber_more_ptr_hwtcl      (0),
    .gen3_coeff_14_nxtber_more_hwtcl          ("g3_coeff_14_nxtber_more"),
    .gen3_coeff_14_nxtber_less_ptr_hwtcl      (0),
    .gen3_coeff_14_nxtber_less_hwtcl          ("g3_coeff_14_nxtber_less"),
    .gen3_coeff_14_reqber_hwtcl               (0),
    .gen3_coeff_14_ber_meas_hwtcl             (0),
    .gen3_coeff_15_hwtcl                      (0),
    .gen3_coeff_15_sel_hwtcl                  ("preset_15"),
    .gen3_coeff_15_preset_hint_hwtcl          (0),
    .gen3_coeff_15_nxtber_more_ptr_hwtcl      (0),
    .gen3_coeff_15_nxtber_more_hwtcl          ("g3_coeff_15_nxtber_more"),
    .gen3_coeff_15_nxtber_less_ptr_hwtcl      (0),
    .gen3_coeff_15_nxtber_less_hwtcl          ("g3_coeff_15_nxtber_less"),
    .gen3_coeff_15_reqber_hwtcl               (0),
    .gen3_coeff_15_ber_meas_hwtcl             (0),
    .gen3_coeff_16_hwtcl                      (0),
    .gen3_coeff_16_sel_hwtcl                  ("preset_16"),
    .gen3_coeff_16_preset_hint_hwtcl          (0),
    .gen3_coeff_16_nxtber_more_ptr_hwtcl      (0),
    .gen3_coeff_16_nxtber_more_hwtcl          ("g3_coeff_16_nxtber_more"),
    .gen3_coeff_16_nxtber_less_ptr_hwtcl      (0),
    .gen3_coeff_16_nxtber_less_hwtcl          ("g3_coeff_16_nxtber_less"),
    .gen3_coeff_16_reqber_hwtcl               (0),
    .gen3_coeff_16_ber_meas_hwtcl             (0),
    .gen3_coeff_17_hwtcl                      (0),
    .gen3_coeff_17_sel_hwtcl                  ("preset_17"),
    .gen3_coeff_17_preset_hint_hwtcl          (0),
    .gen3_coeff_17_nxtber_more_ptr_hwtcl      (0),
    .gen3_coeff_17_nxtber_more_hwtcl          ("g3_coeff_17_nxtber_more"),
    .gen3_coeff_17_nxtber_less_ptr_hwtcl      (0),
    .gen3_coeff_17_nxtber_less_hwtcl          ("g3_coeff_17_nxtber_less"),
    .gen3_coeff_17_reqber_hwtcl               (0),
    .gen3_coeff_17_ber_meas_hwtcl             (0),
    .gen3_coeff_18_hwtcl                      (0),
    .gen3_coeff_18_sel_hwtcl                  ("preset_18"),
    .gen3_coeff_18_preset_hint_hwtcl          (0),
    .gen3_coeff_18_nxtber_more_ptr_hwtcl      (0),
    .gen3_coeff_18_nxtber_more_hwtcl          ("g3_coeff_18_nxtber_more"),
    .gen3_coeff_18_nxtber_less_ptr_hwtcl      (0),
    .gen3_coeff_18_nxtber_less_hwtcl          ("g3_coeff_18_nxtber_less"),
    .gen3_coeff_18_reqber_hwtcl               (0),
    .gen3_coeff_18_ber_meas_hwtcl             (0),
    .gen3_coeff_19_hwtcl                      (0),
    .gen3_coeff_19_sel_hwtcl                  ("preset_19"),
    .gen3_coeff_19_preset_hint_hwtcl          (0),
    .gen3_coeff_19_nxtber_more_ptr_hwtcl      (0),
    .gen3_coeff_19_nxtber_more_hwtcl          ("g3_coeff_19_nxtber_more"),
    .gen3_coeff_19_nxtber_less_ptr_hwtcl      (0),
    .gen3_coeff_19_nxtber_less_hwtcl          ("g3_coeff_19_nxtber_less"),
    .gen3_coeff_19_reqber_hwtcl               (0),
    .gen3_coeff_19_ber_meas_hwtcl             (0),
    .gen3_coeff_20_hwtcl                      (0),
    .gen3_coeff_20_sel_hwtcl                  ("preset_20"),
    .gen3_coeff_20_preset_hint_hwtcl          (0),
    .gen3_coeff_20_nxtber_more_ptr_hwtcl      (0),
    .gen3_coeff_20_nxtber_more_hwtcl          ("g3_coeff_20_nxtber_more"),
    .gen3_coeff_20_nxtber_less_ptr_hwtcl      (0),
    .gen3_coeff_20_nxtber_less_hwtcl          ("g3_coeff_20_nxtber_less"),
    .gen3_coeff_20_reqber_hwtcl               (0),
    .gen3_coeff_20_ber_meas_hwtcl             (0),
    .gen3_coeff_21_hwtcl                      (0),
    .gen3_coeff_21_sel_hwtcl                  ("preset_21"),
    .gen3_coeff_21_preset_hint_hwtcl          (0),
    .gen3_coeff_21_nxtber_more_ptr_hwtcl      (0),
    .gen3_coeff_21_nxtber_more_hwtcl          ("g3_coeff_21_nxtber_more"),
    .gen3_coeff_21_nxtber_less_ptr_hwtcl      (0),
    .gen3_coeff_21_nxtber_less_hwtcl          ("g3_coeff_21_nxtber_less"),
    .gen3_coeff_21_reqber_hwtcl               (0),
    .gen3_coeff_21_ber_meas_hwtcl             (0),
    .gen3_coeff_22_hwtcl                      (0),
    .gen3_coeff_22_sel_hwtcl                  ("preset_22"),
    .gen3_coeff_22_preset_hint_hwtcl          (0),
    .gen3_coeff_22_nxtber_more_ptr_hwtcl      (0),
    .gen3_coeff_22_nxtber_more_hwtcl          ("g3_coeff_22_nxtber_more"),
    .gen3_coeff_22_nxtber_less_ptr_hwtcl      (0),
    .gen3_coeff_22_nxtber_less_hwtcl          ("g3_coeff_22_nxtber_less"),
    .gen3_coeff_22_reqber_hwtcl               (0),
    .gen3_coeff_22_ber_meas_hwtcl             (0),
    .gen3_coeff_23_hwtcl                      (0),
    .gen3_coeff_23_sel_hwtcl                  ("preset_23"),
    .gen3_coeff_23_preset_hint_hwtcl          (0),
    .gen3_coeff_23_nxtber_more_ptr_hwtcl      (0),
    .gen3_coeff_23_nxtber_more_hwtcl          ("g3_coeff_23_nxtber_more"),
    .gen3_coeff_23_nxtber_less_ptr_hwtcl      (0),
    .gen3_coeff_23_nxtber_less_hwtcl          ("g3_coeff_23_nxtber_less"),
    .gen3_coeff_23_reqber_hwtcl               (0),
    .gen3_coeff_23_ber_meas_hwtcl             (0),
    .gen3_coeff_24_hwtcl                      (0),
    .gen3_coeff_24_sel_hwtcl                  ("preset_24"),
    .gen3_coeff_24_preset_hint_hwtcl          (0),
    .gen3_coeff_24_nxtber_more_ptr_hwtcl      (0),
    .gen3_coeff_24_nxtber_more_hwtcl          ("g3_coeff_24_nxtber_more"),
    .gen3_coeff_24_nxtber_less_ptr_hwtcl      (0),
    .gen3_coeff_24_nxtber_less_hwtcl          ("g3_coeff_24_nxtber_less"),
    .gen3_coeff_24_reqber_hwtcl               (0),
    .gen3_coeff_24_ber_meas_hwtcl             (0),
    .hwtcl_override_g3txcoef                  (0),
    .gen3_preset_coeff_1_hwtcl                (0),
    .gen3_preset_coeff_2_hwtcl                (0),
    .gen3_preset_coeff_3_hwtcl                (0),
    .gen3_preset_coeff_4_hwtcl                (0),
    .gen3_preset_coeff_5_hwtcl                (0),
    .gen3_preset_coeff_6_hwtcl                (0),
    .gen3_preset_coeff_7_hwtcl                (0),
    .gen3_preset_coeff_8_hwtcl                (0),
    .gen3_preset_coeff_9_hwtcl                (0),
    .gen3_preset_coeff_10_hwtcl               (0),
    .gen3_preset_coeff_11_hwtcl               (0),
    .gen3_low_freq_hwtcl                      (0),
    .full_swing_hwtcl                         (35),
    .gen3_full_swing_hwtcl                    (35),
    .use_atx_pll_hwtcl                        (0),
    .low_latency_mode_hwtcl                   (0)
  ) dut (
    .npor                   (pcieNPOR_in),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //               npor.npor
    .pin_perst              (pciePERST_in),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //                   .pin_perst
    .lmi_addr               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                lmi.lmi_addr
    .lmi_din                (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .lmi_din
    .lmi_rden               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .lmi_rden
    .lmi_wren               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .lmi_wren
    .lmi_ack                (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .lmi_ack
    .lmi_dout               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .lmi_dout
    .hpg_ctrler             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //          config_tl.hpg_ctrler
    .tl_cfg_add             (tl_cfg_add),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //                   .tl_cfg_add
    .tl_cfg_ctl             (tl_cfg_ctl),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //                   .tl_cfg_ctl
    .tl_cfg_sts             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .tl_cfg_sts
    .cpl_err                (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .cpl_err
    .cpl_pending            (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                   .cpl_pending
    .pm_auxpwr              (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         power_mngt.pm_auxpwr
    .pm_data                (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .pm_data
    .pme_to_cr              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .pme_to_cr
    .pm_event               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .pm_event
    .pme_to_sr              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .pme_to_sr
    .rx_st_sop              (fiData[64]),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //              rx_st.startofpacket
    .rx_st_eop              (fiData[65]),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //                   .endofpacket
    .rx_st_err              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .error
    .rx_st_valid            (fiValid),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                   .valid
    .rx_st_ready            (foReady),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                   .ready
    .rx_st_data             (fiData[63:0]),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //                   .data
    .rx_st_bar              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //          rx_bar_be.rx_st_bar
    .rx_st_be               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .rx_st_be
    .rx_st_mask             (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                   .rx_st_mask
    .tx_st_sop              (txSOP_in),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //              tx_st.startofpacket
    .tx_st_eop              (txEOP_in),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                   .endofpacket
    .tx_st_err              (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                   .error
    .tx_st_valid            (txValid_in),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //                   .valid
    .tx_st_ready            (txReady_out),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                   .ready
    .tx_st_data             (txData_in),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //                   .data
    .tx_cred_datafccp       (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //            tx_cred.tx_cred_datafccp
    .tx_cred_datafcnp       (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .tx_cred_datafcnp
    .tx_cred_datafcp        (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .tx_cred_datafcp
    .tx_cred_fchipcons      (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .tx_cred_fchipcons
    .tx_cred_fcinfinite     (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .tx_cred_fcinfinite
    .tx_cred_hdrfccp        (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .tx_cred_hdrfccp
    .tx_cred_hdrfcnp        (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .tx_cred_hdrfcnp
    .tx_cred_hdrfcp         (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .tx_cred_hdrfcp
    .pld_clk                (pcieClk),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //            pld_clk.clk
    .coreclkout_hip         (pcieClk),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //     coreclkout_hip.clk
    .refclk                 (pcieRefClk_in),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //             refclk.clk
    .reset_status           (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //            hip_rst.reset_status
    .serdes_pll_locked      (pllLocked),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //                   .serdes_pll_locked
    .pld_clk_inuse          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .pld_clk_inuse
    .pld_core_ready         (pllLocked),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //                   .pld_core_ready
    .testin_zero            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .testin_zero
    .reconfig_to_xcvr       (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //   reconfig_to_xcvr.reconfig_to_xcvr
    .reconfig_from_xcvr     (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                // reconfig_from_xcvr.reconfig_from_xcvr
    .rx_in0                 (pcieRX_in[0]),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //         hip_serial.rx_in0
    .rx_in1                 (pcieRX_in[1]),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //                   .rx_in1
    .rx_in2                 (pcieRX_in[2]),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //                   .rx_in2
    .rx_in3                 (pcieRX_in[3]),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //                   .rx_in3
    .tx_out0                (pcieTX_out[0]),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //                   .tx_out0
    .tx_out1                (pcieTX_out[1]),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //                   .tx_out1
    .tx_out2                (pcieTX_out[2]),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //                   .tx_out2
    .tx_out3                (pcieTX_out[3]),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //                   .tx_out3
    .sim_pipe_pclk_in       (hip_pipe_sim_pipe_pclk_in),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //           hip_pipe.sim_pipe_pclk_in
    .sim_pipe_rate          (hip_pipe_sim_pipe_rate),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //                   .sim_pipe_rate
    .sim_ltssmstate         (hip_pipe_sim_ltssmstate),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                   .sim_ltssmstate
    .eidleinfersel0         (hip_pipe_eidleinfersel0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                   .eidleinfersel0
    .eidleinfersel1         (hip_pipe_eidleinfersel1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                   .eidleinfersel1
    .eidleinfersel2         (hip_pipe_eidleinfersel2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                   .eidleinfersel2
    .eidleinfersel3         (hip_pipe_eidleinfersel3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                   .eidleinfersel3
    .powerdown0             (hip_pipe_powerdown0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                   .powerdown0
    .powerdown1             (hip_pipe_powerdown1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                   .powerdown1
    .powerdown2             (hip_pipe_powerdown2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                   .powerdown2
    .powerdown3             (hip_pipe_powerdown3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                   .powerdown3
    .rxpolarity0            (hip_pipe_rxpolarity0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                   .rxpolarity0
    .rxpolarity1            (hip_pipe_rxpolarity1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                   .rxpolarity1
    .rxpolarity2            (hip_pipe_rxpolarity2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                   .rxpolarity2
    .rxpolarity3            (hip_pipe_rxpolarity3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                   .rxpolarity3
    .txcompl0               (hip_pipe_txcompl0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .txcompl0
    .txcompl1               (hip_pipe_txcompl1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .txcompl1
    .txcompl2               (hip_pipe_txcompl2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .txcompl2
    .txcompl3               (hip_pipe_txcompl3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .txcompl3
    .txdata0                (hip_pipe_txdata0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .txdata0
    .txdata1                (hip_pipe_txdata1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .txdata1
    .txdata2                (hip_pipe_txdata2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .txdata2
    .txdata3                (hip_pipe_txdata3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .txdata3
    .txdatak0               (hip_pipe_txdatak0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .txdatak0
    .txdatak1               (hip_pipe_txdatak1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .txdatak1
    .txdatak2               (hip_pipe_txdatak2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .txdatak2
    .txdatak3               (hip_pipe_txdatak3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .txdatak3
    .txdetectrx0            (hip_pipe_txdetectrx0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                   .txdetectrx0
    .txdetectrx1            (hip_pipe_txdetectrx1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                   .txdetectrx1
    .txdetectrx2            (hip_pipe_txdetectrx2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                   .txdetectrx2
    .txdetectrx3            (hip_pipe_txdetectrx3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                   .txdetectrx3
    .txelecidle0            (hip_pipe_txelecidle0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                   .txelecidle0
    .txelecidle1            (hip_pipe_txelecidle1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                   .txelecidle1
    .txelecidle2            (hip_pipe_txelecidle2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                   .txelecidle2
    .txelecidle3            (hip_pipe_txelecidle3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                   .txelecidle3
    .txdeemph0              (hip_pipe_txdeemph0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                   .txdeemph0
    .txdeemph1              (hip_pipe_txdeemph1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                   .txdeemph1
    .txdeemph2              (hip_pipe_txdeemph2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                   .txdeemph2
    .txdeemph3              (hip_pipe_txdeemph3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                   .txdeemph3
    .txmargin0              (hip_pipe_txmargin0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                   .txmargin0
    .txmargin1              (hip_pipe_txmargin1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                   .txmargin1
    .txmargin2              (hip_pipe_txmargin2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                   .txmargin2
    .txmargin3              (hip_pipe_txmargin3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                   .txmargin3
    .txswing0               (hip_pipe_txswing0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .txswing0
    .txswing1               (hip_pipe_txswing1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .txswing1
    .txswing2               (hip_pipe_txswing2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .txswing2
    .txswing3               (hip_pipe_txswing3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .txswing3
    .phystatus0             (hip_pipe_phystatus0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                   .phystatus0
    .phystatus1             (hip_pipe_phystatus1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                   .phystatus1
    .phystatus2             (hip_pipe_phystatus2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                   .phystatus2
    .phystatus3             (hip_pipe_phystatus3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                   .phystatus3
    .rxdata0                (hip_pipe_rxdata0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .rxdata0
    .rxdata1                (hip_pipe_rxdata1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .rxdata1
    .rxdata2                (hip_pipe_rxdata2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .rxdata2
    .rxdata3                (hip_pipe_rxdata3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .rxdata3
    .rxdatak0               (hip_pipe_rxdatak0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .rxdatak0
    .rxdatak1               (hip_pipe_rxdatak1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .rxdatak1
    .rxdatak2               (hip_pipe_rxdatak2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .rxdatak2
    .rxdatak3               (hip_pipe_rxdatak3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .rxdatak3
    .rxelecidle0            (hip_pipe_rxelecidle0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                   .rxelecidle0
    .rxelecidle1            (hip_pipe_rxelecidle1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                   .rxelecidle1
    .rxelecidle2            (hip_pipe_rxelecidle2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                   .rxelecidle2
    .rxelecidle3            (hip_pipe_rxelecidle3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                   .rxelecidle3
    .rxstatus0              (hip_pipe_rxstatus0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                   .rxstatus0
    .rxstatus1              (hip_pipe_rxstatus1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                   .rxstatus1
    .rxstatus2              (hip_pipe_rxstatus2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                   .rxstatus2
    .rxstatus3              (hip_pipe_rxstatus3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                   .rxstatus3
    .rxvalid0               (hip_pipe_rxvalid0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .rxvalid0
    .rxvalid1               (hip_pipe_rxvalid1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .rxvalid1
    .rxvalid2               (hip_pipe_rxvalid2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .rxvalid2
    .rxvalid3               (hip_pipe_rxvalid3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .rxvalid3
    .app_int_sts            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //            int_msi.app_int_sts
    .app_msi_num            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .app_msi_num
    .app_msi_req            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .app_msi_req
    .app_msi_tc             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .app_msi_tc
    .app_int_ack            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .app_int_ack
    .app_msi_ack            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .app_msi_ack
    .test_in                (hip_ctrl_test_in),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //           hip_ctrl.test_in
    .simu_mode_pipe         (hip_ctrl_simu_mode_pipe),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                   .simu_mode_pipe
    .derr_cor_ext_rcv       (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         hip_status.derr_cor_ext_rcv
    .derr_cor_ext_rpl       (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .derr_cor_ext_rpl
    .derr_rpl               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .derr_rpl
    .dlup                   (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .dlup
    .dlup_exit              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .dlup_exit
    .ev128ns                (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .ev128ns
    .ev1us                  (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .ev1us
    .hotrst_exit            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .hotrst_exit
    .int_status             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .int_status
    .l2_exit                (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .l2_exit
    .lane_act               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .lane_act
    .ltssmstate             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .ltssmstate
    .rx_par_err             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .rx_par_err
    .tx_par_err             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .tx_par_err
    .cfg_par_err            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .cfg_par_err
    .ko_cpl_spc_header      (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .ko_cpl_spc_header
    .ko_cpl_spc_data        (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .ko_cpl_spc_data
    .currentspeed           (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //   hip_currentspeed.currentspeed
    .rx_st_empty            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .rx_st_parity           (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .tx_st_empty            (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //        (terminated)
    .tx_st_parity           (8'b00000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //        (terminated)
    .tx_cons_cred_sel       (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .sim_pipe_pclk_out      (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .rx_in4                 (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .rx_in5                 (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .rx_in6                 (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .rx_in7                 (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .tx_out4                (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .tx_out5                (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .tx_out6                (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .tx_out7                (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .eidleinfersel4         (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .eidleinfersel5         (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .eidleinfersel6         (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .eidleinfersel7         (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .powerdown4             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .powerdown5             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .powerdown6             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .powerdown7             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .rxpolarity4            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .rxpolarity5            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .rxpolarity6            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .rxpolarity7            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .txcompl4               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .txcompl5               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .txcompl6               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .txcompl7               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .txdata4                (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .txdata5                (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .txdata6                (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .txdata7                (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .txdatak4               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .txdatak5               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .txdatak6               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .txdatak7               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .txdetectrx4            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .txdetectrx5            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .txdetectrx6            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .txdetectrx7            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .txelecidle4            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .txelecidle5            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .txelecidle6            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .txelecidle7            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .txdeemph4              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .txdeemph5              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .txdeemph6              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .txdeemph7              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .txmargin4              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .txmargin5              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .txmargin6              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .txmargin7              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .txswing4               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .txswing5               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .txswing6               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .txswing7               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .phystatus4             (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .phystatus5             (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .phystatus6             (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .phystatus7             (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .rxdata4                (8'b00000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //        (terminated)
    .rxdata5                (8'b00000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //        (terminated)
    .rxdata6                (8'b00000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //        (terminated)
    .rxdata7                (8'b00000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //        (terminated)
    .rxdatak4               (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .rxdatak5               (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .rxdatak6               (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .rxdatak7               (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .rxelecidle4            (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .rxelecidle5            (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .rxelecidle6            (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .rxelecidle7            (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .rxstatus4              (3'b000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //        (terminated)
    .rxstatus5              (3'b000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //        (terminated)
    .rxstatus6              (3'b000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //        (terminated)
    .rxstatus7              (3'b000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //        (terminated)
    .rxvalid4               (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .rxvalid5               (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .rxvalid6               (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .rxvalid7               (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .rxdataskip0            (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .rxdataskip1            (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .rxdataskip2            (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .rxdataskip3            (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .rxdataskip4            (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .rxdataskip5            (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .rxdataskip6            (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .rxdataskip7            (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .rxblkst0               (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .rxblkst1               (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .rxblkst2               (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .rxblkst3               (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .rxblkst4               (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .rxblkst5               (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .rxblkst6               (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .rxblkst7               (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .rxsynchd0              (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //        (terminated)
    .rxsynchd1              (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //        (terminated)
    .rxsynchd2              (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //        (terminated)
    .rxsynchd3              (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //        (terminated)
    .rxsynchd4              (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //        (terminated)
    .rxsynchd5              (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //        (terminated)
    .rxsynchd6              (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //        (terminated)
    .rxsynchd7              (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //        (terminated)
    .rxfreqlocked0          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .rxfreqlocked1          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .rxfreqlocked2          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .rxfreqlocked3          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .rxfreqlocked4          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .rxfreqlocked5          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .rxfreqlocked6          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .rxfreqlocked7          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .currentcoeff0          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .currentcoeff1          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .currentcoeff2          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .currentcoeff3          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .currentcoeff4          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .currentcoeff5          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .currentcoeff6          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .currentcoeff7          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .currentrxpreset0       (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .currentrxpreset1       (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .currentrxpreset2       (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .currentrxpreset3       (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .currentrxpreset4       (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .currentrxpreset5       (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .currentrxpreset6       (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .currentrxpreset7       (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .txsynchd0              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .txsynchd1              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .txsynchd2              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .txsynchd3              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .txsynchd4              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .txsynchd5              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .txsynchd6              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .txsynchd7              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .txblkst0               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .txblkst1               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .txblkst2               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .txblkst3               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .txblkst4               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .txblkst5               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .txblkst6               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .txblkst7               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .aer_msi_num            (5'b00000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //        (terminated)
    .pex_msi_num            (5'b00000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //        (terminated)
    .serr_out               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .hip_reconfig_clk       (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .hip_reconfig_rst_n     (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .hip_reconfig_address   (10'b0000000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //        (terminated)
    .hip_reconfig_read      (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .hip_reconfig_write     (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .hip_reconfig_writedata (16'b0000000000000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .hip_reconfig_byte_en   (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //        (terminated)
    .ser_shift_load         (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .interface_sel          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .cfgbp_link2csr         (13'b0000000000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //        (terminated)
    .cfgbp_comclk_reg       (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .cfgbp_extsy_reg        (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .cfgbp_max_pload        (3'b000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //        (terminated)
    .cfgbp_tx_ecrcgen       (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .cfgbp_rx_ecrchk        (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .cfgbp_secbus           (8'b00000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //        (terminated)
    .cfgbp_linkcsr_bit0     (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .cfgbp_tx_req_pm        (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .cfgbp_tx_typ_pm        (3'b000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //        (terminated)
    .cfgbp_req_phypm        (4'b0000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //        (terminated)
    .cfgbp_req_phycfg       (4'b0000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //        (terminated)
    .cfgbp_vc0_tcmap_pld    (7'b0000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //        (terminated)
    .cfgbp_inh_dllp         (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .cfgbp_inh_tx_tlp       (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .cfgbp_req_wake         (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .cfgbp_link3_ctl        (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //        (terminated)
    .cseb_rddata            (32'b00000000000000000000000000000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .cseb_rdresponse        (5'b00000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //        (terminated)
    .cseb_waitrequest       (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .cseb_wrresponse        (5'b00000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //        (terminated)
    .cseb_wrresp_valid      (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .cseb_rddata_parity     (4'b0000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //        (terminated)
    .reservedin             (32'b00000000000000000000000000000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
    .tlbfm_in               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
    .tlbfm_out              (1001'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000), //        (terminated)
    .rxfc_cplbuf_ovf        ()                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //        (terminated)
  );

endmodule
