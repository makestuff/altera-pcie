//
// Copyright (C) 2014, 2017-2018 Chris McClelland
//
// Permission is hereby granted, free of charge, to any person obtaining a copy of this software
// and associated documentation files (the "Software"), to deal in the Software without
// restriction, including without limitation the rights to use, copy, modify, merge, publish,
// distribute, sublicense, and/or sell copies of the Software, and to permit persons to whom the
// Software is furnished to do so, subject to the following conditions:
//
// The above copyright  notice and this permission notice  shall be included in all copies or
// substantial portions of the Software.
//
// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR IMPLIED, INCLUDING
// BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND
// NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM,
// DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE SOFTWARE.
//
`timescale 1 ps / 1 ps
module pcie_sv_tb;

  wire  [31:0] dut_pcie_tb_hip_ctrl_test_in;          // DUT_pcie_tb:test_in -> pcie_sv_inst:hip_ctrl_test_in
  wire         dut_pcie_tb_hip_ctrl_simu_mode_pipe;   // DUT_pcie_tb:simu_mode_pipe -> pcie_sv_inst:hip_ctrl_simu_mode_pipe
  wire   [7:0] pcie_sv_inst_hip_pipe_txdata3;         // pcie_sv_inst:hip_pipe_txdata3 -> DUT_pcie_tb:txdata3
  wire   [7:0] pcie_sv_inst_hip_pipe_txdata2;         // pcie_sv_inst:hip_pipe_txdata2 -> DUT_pcie_tb:txdata2
  wire   [7:0] pcie_sv_inst_hip_pipe_txdata1;         // pcie_sv_inst:hip_pipe_txdata1 -> DUT_pcie_tb:txdata1
  wire   [7:0] pcie_sv_inst_hip_pipe_txdata0;         // pcie_sv_inst:hip_pipe_txdata0 -> DUT_pcie_tb:txdata0
  wire   [2:0] dut_pcie_tb_hip_pipe_rxstatus2;        // DUT_pcie_tb:rxstatus2 -> pcie_sv_inst:hip_pipe_rxstatus2
  wire   [2:0] dut_pcie_tb_hip_pipe_rxstatus3;        // DUT_pcie_tb:rxstatus3 -> pcie_sv_inst:hip_pipe_rxstatus3
  wire         pcie_sv_inst_hip_pipe_rxpolarity2;     // pcie_sv_inst:hip_pipe_rxpolarity2 -> DUT_pcie_tb:rxpolarity2
  wire   [2:0] dut_pcie_tb_hip_pipe_rxstatus0;        // DUT_pcie_tb:rxstatus0 -> pcie_sv_inst:hip_pipe_rxstatus0
  wire         pcie_sv_inst_hip_pipe_rxpolarity3;     // pcie_sv_inst:hip_pipe_rxpolarity3 -> DUT_pcie_tb:rxpolarity3
  wire         dut_pcie_tb_hip_pipe_rxelecidle3;      // DUT_pcie_tb:rxelecidle3 -> pcie_sv_inst:hip_pipe_rxelecidle3
  wire   [2:0] dut_pcie_tb_hip_pipe_rxstatus1;        // DUT_pcie_tb:rxstatus1 -> pcie_sv_inst:hip_pipe_rxstatus1
  wire         pcie_sv_inst_hip_pipe_rxpolarity0;     // pcie_sv_inst:hip_pipe_rxpolarity0 -> DUT_pcie_tb:rxpolarity0
  wire         dut_pcie_tb_hip_pipe_rxelecidle2;      // DUT_pcie_tb:rxelecidle2 -> pcie_sv_inst:hip_pipe_rxelecidle2
  wire         pcie_sv_inst_hip_pipe_rxpolarity1;     // pcie_sv_inst:hip_pipe_rxpolarity1 -> DUT_pcie_tb:rxpolarity1
  wire         dut_pcie_tb_hip_pipe_rxelecidle1;      // DUT_pcie_tb:rxelecidle1 -> pcie_sv_inst:hip_pipe_rxelecidle1
  wire         dut_pcie_tb_hip_pipe_rxelecidle0;      // DUT_pcie_tb:rxelecidle0 -> pcie_sv_inst:hip_pipe_rxelecidle0
  wire         dut_pcie_tb_hip_pipe_phystatus0;       // DUT_pcie_tb:phystatus0 -> pcie_sv_inst:hip_pipe_phystatus0
  wire         pcie_sv_inst_hip_pipe_txswing3;        // pcie_sv_inst:hip_pipe_txswing3 -> DUT_pcie_tb:txswing3
  wire         dut_pcie_tb_hip_pipe_phystatus1;       // DUT_pcie_tb:phystatus1 -> pcie_sv_inst:hip_pipe_phystatus1
  wire         pcie_sv_inst_hip_pipe_txswing2;        // pcie_sv_inst:hip_pipe_txswing2 -> DUT_pcie_tb:txswing2
  wire         dut_pcie_tb_hip_pipe_phystatus2;       // DUT_pcie_tb:phystatus2 -> pcie_sv_inst:hip_pipe_phystatus2
  wire         pcie_sv_inst_hip_pipe_txswing1;        // pcie_sv_inst:hip_pipe_txswing1 -> DUT_pcie_tb:txswing1
  wire         pcie_sv_inst_hip_pipe_txswing0;        // pcie_sv_inst:hip_pipe_txswing0 -> DUT_pcie_tb:txswing0
  wire         pcie_sv_inst_hip_pipe_txcompl0;        // pcie_sv_inst:hip_pipe_txcompl0 -> DUT_pcie_tb:txcompl0
  wire         dut_pcie_tb_hip_pipe_phystatus3;       // DUT_pcie_tb:phystatus3 -> pcie_sv_inst:hip_pipe_phystatus3
  wire         pcie_sv_inst_hip_pipe_txcompl3;        // pcie_sv_inst:hip_pipe_txcompl3 -> DUT_pcie_tb:txcompl3
  wire         pcie_sv_inst_hip_pipe_txcompl2;        // pcie_sv_inst:hip_pipe_txcompl2 -> DUT_pcie_tb:txcompl2
  wire         pcie_sv_inst_hip_pipe_txcompl1;        // pcie_sv_inst:hip_pipe_txcompl1 -> DUT_pcie_tb:txcompl1
  wire   [2:0] pcie_sv_inst_hip_pipe_txmargin1;       // pcie_sv_inst:hip_pipe_txmargin1 -> DUT_pcie_tb:txmargin1
  wire   [2:0] pcie_sv_inst_hip_pipe_txmargin0;       // pcie_sv_inst:hip_pipe_txmargin0 -> DUT_pcie_tb:txmargin0
  wire   [2:0] pcie_sv_inst_hip_pipe_eidleinfersel1;  // pcie_sv_inst:hip_pipe_eidleinfersel1 -> DUT_pcie_tb:eidleinfersel1
  wire   [2:0] pcie_sv_inst_hip_pipe_eidleinfersel2;  // pcie_sv_inst:hip_pipe_eidleinfersel2 -> DUT_pcie_tb:eidleinfersel2
  wire         pcie_sv_inst_hip_pipe_txdeemph0;       // pcie_sv_inst:hip_pipe_txdeemph0 -> DUT_pcie_tb:txdeemph0
  wire   [2:0] pcie_sv_inst_hip_pipe_eidleinfersel3;  // pcie_sv_inst:hip_pipe_eidleinfersel3 -> DUT_pcie_tb:eidleinfersel3
  wire         pcie_sv_inst_hip_pipe_txdeemph3;       // pcie_sv_inst:hip_pipe_txdeemph3 -> DUT_pcie_tb:txdeemph3
  wire         pcie_sv_inst_hip_pipe_txdeemph1;       // pcie_sv_inst:hip_pipe_txdeemph1 -> DUT_pcie_tb:txdeemph1
  wire   [2:0] pcie_sv_inst_hip_pipe_eidleinfersel0;  // pcie_sv_inst:hip_pipe_eidleinfersel0 -> DUT_pcie_tb:eidleinfersel0
  wire         pcie_sv_inst_hip_pipe_txdeemph2;       // pcie_sv_inst:hip_pipe_txdeemph2 -> DUT_pcie_tb:txdeemph2
  wire   [7:0] dut_pcie_tb_hip_pipe_rxdata2;          // DUT_pcie_tb:rxdata2 -> pcie_sv_inst:hip_pipe_rxdata2
  wire   [7:0] dut_pcie_tb_hip_pipe_rxdata3;          // DUT_pcie_tb:rxdata3 -> pcie_sv_inst:hip_pipe_rxdata3
  wire   [7:0] dut_pcie_tb_hip_pipe_rxdata0;          // DUT_pcie_tb:rxdata0 -> pcie_sv_inst:hip_pipe_rxdata0
  wire         pcie_sv_inst_hip_pipe_txelecidle0;     // pcie_sv_inst:hip_pipe_txelecidle0 -> DUT_pcie_tb:txelecidle0
  wire   [7:0] dut_pcie_tb_hip_pipe_rxdata1;          // DUT_pcie_tb:rxdata1 -> pcie_sv_inst:hip_pipe_rxdata1
  wire         pcie_sv_inst_hip_pipe_txelecidle1;     // pcie_sv_inst:hip_pipe_txelecidle1 -> DUT_pcie_tb:txelecidle1
  wire         pcie_sv_inst_hip_pipe_txelecidle2;     // pcie_sv_inst:hip_pipe_txelecidle2 -> DUT_pcie_tb:txelecidle2
  wire         dut_pcie_tb_hip_pipe_sim_pipe_pclk_in; // DUT_pcie_tb:sim_pipe_pclk_in -> pcie_sv_inst:hip_pipe_sim_pipe_pclk_in
  wire         pcie_sv_inst_hip_pipe_txelecidle3;     // pcie_sv_inst:hip_pipe_txelecidle3 -> DUT_pcie_tb:txelecidle3
  wire   [1:0] pcie_sv_inst_hip_pipe_sim_pipe_rate;   // pcie_sv_inst:hip_pipe_sim_pipe_rate -> DUT_pcie_tb:sim_pipe_rate
  wire         pcie_sv_inst_hip_pipe_txdetectrx2;     // pcie_sv_inst:hip_pipe_txdetectrx2 -> DUT_pcie_tb:txdetectrx2
  wire         pcie_sv_inst_hip_pipe_txdetectrx1;     // pcie_sv_inst:hip_pipe_txdetectrx1 -> DUT_pcie_tb:txdetectrx1
  wire   [2:0] pcie_sv_inst_hip_pipe_txmargin3;       // pcie_sv_inst:hip_pipe_txmargin3 -> DUT_pcie_tb:txmargin3
  wire         pcie_sv_inst_hip_pipe_txdetectrx3;     // pcie_sv_inst:hip_pipe_txdetectrx3 -> DUT_pcie_tb:txdetectrx3
  wire   [2:0] pcie_sv_inst_hip_pipe_txmargin2;       // pcie_sv_inst:hip_pipe_txmargin2 -> DUT_pcie_tb:txmargin2
  wire         pcie_sv_inst_hip_pipe_txdetectrx0;     // pcie_sv_inst:hip_pipe_txdetectrx0 -> DUT_pcie_tb:txdetectrx0
  wire   [1:0] pcie_sv_inst_hip_pipe_powerdown3;      // pcie_sv_inst:hip_pipe_powerdown3 -> DUT_pcie_tb:powerdown3
  wire   [1:0] pcie_sv_inst_hip_pipe_powerdown0;      // pcie_sv_inst:hip_pipe_powerdown0 -> DUT_pcie_tb:powerdown0
  wire   [1:0] pcie_sv_inst_hip_pipe_powerdown1;      // pcie_sv_inst:hip_pipe_powerdown1 -> DUT_pcie_tb:powerdown1
  wire   [1:0] pcie_sv_inst_hip_pipe_powerdown2;      // pcie_sv_inst:hip_pipe_powerdown2 -> DUT_pcie_tb:powerdown2
  wire   [4:0] pcie_sv_inst_hip_pipe_sim_ltssmstate;  // pcie_sv_inst:hip_pipe_sim_ltssmstate -> DUT_pcie_tb:sim_ltssmstate
  wire         dut_pcie_tb_hip_pipe_rxvalid3;         // DUT_pcie_tb:rxvalid3 -> pcie_sv_inst:hip_pipe_rxvalid3
  wire         dut_pcie_tb_hip_pipe_rxvalid2;         // DUT_pcie_tb:rxvalid2 -> pcie_sv_inst:hip_pipe_rxvalid2
  wire         dut_pcie_tb_hip_pipe_rxvalid1;         // DUT_pcie_tb:rxvalid1 -> pcie_sv_inst:hip_pipe_rxvalid1
  wire         dut_pcie_tb_hip_pipe_rxvalid0;         // DUT_pcie_tb:rxvalid0 -> pcie_sv_inst:hip_pipe_rxvalid0
  wire         pcie_sv_inst_hip_pipe_txdatak2;        // pcie_sv_inst:hip_pipe_txdatak2 -> DUT_pcie_tb:txdatak2
  wire         pcie_sv_inst_hip_pipe_txdatak1;        // pcie_sv_inst:hip_pipe_txdatak1 -> DUT_pcie_tb:txdatak1
  wire         pcie_sv_inst_hip_pipe_txdatak3;        // pcie_sv_inst:hip_pipe_txdatak3 -> DUT_pcie_tb:txdatak3
  wire         dut_pcie_tb_hip_pipe_rxdatak2;         // DUT_pcie_tb:rxdatak2 -> pcie_sv_inst:hip_pipe_rxdatak2
  wire         dut_pcie_tb_hip_pipe_rxdatak1;         // DUT_pcie_tb:rxdatak1 -> pcie_sv_inst:hip_pipe_rxdatak1
  wire         pcie_sv_inst_hip_pipe_txdatak0;        // pcie_sv_inst:hip_pipe_txdatak0 -> DUT_pcie_tb:txdatak0
  wire         dut_pcie_tb_hip_pipe_rxdatak0;         // DUT_pcie_tb:rxdatak0 -> pcie_sv_inst:hip_pipe_rxdatak0
  wire         dut_pcie_tb_hip_pipe_rxdatak3;         // DUT_pcie_tb:rxdatak3 -> pcie_sv_inst:hip_pipe_rxdatak3

  // External signals
  logic pcieRefClk;
  logic pcieNPOR;
  logic pciePERST;

  // Application interface
  logic        pcieClk;    // 125MHz core clock from PCIe PLL
  logic[12:0]  cfgBusDev;  // the device ID assigned to the FPGA on enumeration

  logic[63:0]  rxData;     // incoming requests from the CPU
  logic        rxSOP;
  logic        rxEOP;
  logic        rxValid;
  logic        rxReady;

  logic[63:0]  txData;     // outgoing responses from the FPGA
  logic        txSOP;
  logic        txEOP;
  logic        txValid;
  logic        txReady;

  // The thing which actually drives the bus from the FPGA side
  pcie_app pcie_app (
    .pcieClk_in    (pcieClk),
    .cfgBusDev_in  (cfgBusDev),

    .rxData_in     (rxData),
    .rxValid_in    (rxValid),
    .rxReady_out   (rxReady),
    .rxSOP_in      (rxSOP),
    .rxEOP_in      (rxEOP),

    .txData_out    (txData),
    .txValid_out   (txValid),
    .txReady_in    (txReady),
    .txSOP_out     (txSOP),
    .txEOP_out     (txEOP)
  );

  // Testbench which simulates the behaviour of a Root-Port (i.e a host PC). Ultimately, this
  // executes the bus activity specified in altpcietb_bfm_driver_chaining.v.
  altpcie_tbed_sv_hwtcl #(
    .lane_mask_hwtcl                      ("x4"),
    .gen123_lane_rate_mode_hwtcl          ("Gen1 (2.5 Gbps)"),
    .port_type_hwtcl                      ("Native endpoint"),
    .pll_refclk_freq_hwtcl                ("100 MHz"),
    .apps_type_hwtcl                      (2),
    .serial_sim_hwtcl                     (0),
    .enable_pipe32_sim_hwtcl              (0),
    .enable_tl_only_sim_hwtcl             (0),
    .deemphasis_enable_hwtcl              ("false"),
    .pld_clk_MHz                          (1250),
    .millisecond_cycle_count_hwtcl        (124250),
    .use_crc_forwarding_hwtcl             (0),
    .ecrc_check_capable_hwtcl             (0),
    .ecrc_gen_capable_hwtcl               (0),
    .enable_pipe32_phyip_ser_driver_hwtcl (0)
  ) dut_pcie_tb (
    .npor             (pcieNPOR),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //       npor.npor
    .pin_perst        (pciePERST),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //           .pin_perst
    .refclk           (pcieRefClk),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //     refclk.clk
    .sim_pipe_pclk_in (dut_pcie_tb_hip_pipe_sim_pipe_pclk_in),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //   hip_pipe.sim_pipe_pclk_in
    .sim_pipe_rate    (pcie_sv_inst_hip_pipe_sim_pipe_rate),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //           .sim_pipe_rate
    .sim_ltssmstate   (pcie_sv_inst_hip_pipe_sim_ltssmstate),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //           .sim_ltssmstate
    .eidleinfersel0   (pcie_sv_inst_hip_pipe_eidleinfersel0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //           .eidleinfersel0
    .eidleinfersel1   (pcie_sv_inst_hip_pipe_eidleinfersel1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //           .eidleinfersel1
    .eidleinfersel2   (pcie_sv_inst_hip_pipe_eidleinfersel2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //           .eidleinfersel2
    .eidleinfersel3   (pcie_sv_inst_hip_pipe_eidleinfersel3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //           .eidleinfersel3
    .powerdown0       (pcie_sv_inst_hip_pipe_powerdown0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //           .powerdown0
    .powerdown1       (pcie_sv_inst_hip_pipe_powerdown1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //           .powerdown1
    .powerdown2       (pcie_sv_inst_hip_pipe_powerdown2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //           .powerdown2
    .powerdown3       (pcie_sv_inst_hip_pipe_powerdown3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //           .powerdown3
    .rxpolarity0      (pcie_sv_inst_hip_pipe_rxpolarity0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //           .rxpolarity0
    .rxpolarity1      (pcie_sv_inst_hip_pipe_rxpolarity1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //           .rxpolarity1
    .rxpolarity2      (pcie_sv_inst_hip_pipe_rxpolarity2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //           .rxpolarity2
    .rxpolarity3      (pcie_sv_inst_hip_pipe_rxpolarity3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //           .rxpolarity3
    .txcompl0         (pcie_sv_inst_hip_pipe_txcompl0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //           .txcompl0
    .txcompl1         (pcie_sv_inst_hip_pipe_txcompl1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //           .txcompl1
    .txcompl2         (pcie_sv_inst_hip_pipe_txcompl2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //           .txcompl2
    .txcompl3         (pcie_sv_inst_hip_pipe_txcompl3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //           .txcompl3
    .txdata0          (pcie_sv_inst_hip_pipe_txdata0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //           .txdata0
    .txdata1          (pcie_sv_inst_hip_pipe_txdata1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //           .txdata1
    .txdata2          (pcie_sv_inst_hip_pipe_txdata2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //           .txdata2
    .txdata3          (pcie_sv_inst_hip_pipe_txdata3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //           .txdata3
    .txdatak0         (pcie_sv_inst_hip_pipe_txdatak0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //           .txdatak0
    .txdatak1         (pcie_sv_inst_hip_pipe_txdatak1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //           .txdatak1
    .txdatak2         (pcie_sv_inst_hip_pipe_txdatak2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //           .txdatak2
    .txdatak3         (pcie_sv_inst_hip_pipe_txdatak3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //           .txdatak3
    .txdetectrx0      (pcie_sv_inst_hip_pipe_txdetectrx0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //           .txdetectrx0
    .txdetectrx1      (pcie_sv_inst_hip_pipe_txdetectrx1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //           .txdetectrx1
    .txdetectrx2      (pcie_sv_inst_hip_pipe_txdetectrx2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //           .txdetectrx2
    .txdetectrx3      (pcie_sv_inst_hip_pipe_txdetectrx3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //           .txdetectrx3
    .txelecidle0      (pcie_sv_inst_hip_pipe_txelecidle0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //           .txelecidle0
    .txelecidle1      (pcie_sv_inst_hip_pipe_txelecidle1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //           .txelecidle1
    .txelecidle2      (pcie_sv_inst_hip_pipe_txelecidle2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //           .txelecidle2
    .txelecidle3      (pcie_sv_inst_hip_pipe_txelecidle3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //           .txelecidle3
    .txdeemph0        (pcie_sv_inst_hip_pipe_txdeemph0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //           .txdeemph0
    .txdeemph1        (pcie_sv_inst_hip_pipe_txdeemph1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //           .txdeemph1
    .txdeemph2        (pcie_sv_inst_hip_pipe_txdeemph2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //           .txdeemph2
    .txdeemph3        (pcie_sv_inst_hip_pipe_txdeemph3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //           .txdeemph3
    .txmargin0        (pcie_sv_inst_hip_pipe_txmargin0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //           .txmargin0
    .txmargin1        (pcie_sv_inst_hip_pipe_txmargin1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //           .txmargin1
    .txmargin2        (pcie_sv_inst_hip_pipe_txmargin2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //           .txmargin2
    .txmargin3        (pcie_sv_inst_hip_pipe_txmargin3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //           .txmargin3
    .txswing0         (pcie_sv_inst_hip_pipe_txswing0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //           .txswing0
    .txswing1         (pcie_sv_inst_hip_pipe_txswing1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //           .txswing1
    .txswing2         (pcie_sv_inst_hip_pipe_txswing2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //           .txswing2
    .txswing3         (pcie_sv_inst_hip_pipe_txswing3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //           .txswing3
    .phystatus0       (dut_pcie_tb_hip_pipe_phystatus0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //           .phystatus0
    .phystatus1       (dut_pcie_tb_hip_pipe_phystatus1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //           .phystatus1
    .phystatus2       (dut_pcie_tb_hip_pipe_phystatus2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //           .phystatus2
    .phystatus3       (dut_pcie_tb_hip_pipe_phystatus3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //           .phystatus3
    .rxdata0          (dut_pcie_tb_hip_pipe_rxdata0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //           .rxdata0
    .rxdata1          (dut_pcie_tb_hip_pipe_rxdata1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //           .rxdata1
    .rxdata2          (dut_pcie_tb_hip_pipe_rxdata2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //           .rxdata2
    .rxdata3          (dut_pcie_tb_hip_pipe_rxdata3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //           .rxdata3
    .rxdatak0         (dut_pcie_tb_hip_pipe_rxdatak0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //           .rxdatak0
    .rxdatak1         (dut_pcie_tb_hip_pipe_rxdatak1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //           .rxdatak1
    .rxdatak2         (dut_pcie_tb_hip_pipe_rxdatak2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //           .rxdatak2
    .rxdatak3         (dut_pcie_tb_hip_pipe_rxdatak3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //           .rxdatak3
    .rxelecidle0      (dut_pcie_tb_hip_pipe_rxelecidle0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //           .rxelecidle0
    .rxelecidle1      (dut_pcie_tb_hip_pipe_rxelecidle1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //           .rxelecidle1
    .rxelecidle2      (dut_pcie_tb_hip_pipe_rxelecidle2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //           .rxelecidle2
    .rxelecidle3      (dut_pcie_tb_hip_pipe_rxelecidle3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //           .rxelecidle3
    .rxstatus0        (dut_pcie_tb_hip_pipe_rxstatus0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //           .rxstatus0
    .rxstatus1        (dut_pcie_tb_hip_pipe_rxstatus1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //           .rxstatus1
    .rxstatus2        (dut_pcie_tb_hip_pipe_rxstatus2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //           .rxstatus2
    .rxstatus3        (dut_pcie_tb_hip_pipe_rxstatus3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //           .rxstatus3
    .rxvalid0         (dut_pcie_tb_hip_pipe_rxvalid0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //           .rxvalid0
    .rxvalid1         (dut_pcie_tb_hip_pipe_rxvalid1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //           .rxvalid1
    .rxvalid2         (dut_pcie_tb_hip_pipe_rxvalid2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //           .rxvalid2
    .rxvalid3         (dut_pcie_tb_hip_pipe_rxvalid3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //           .rxvalid3
    .rx_in0           (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                // hip_serial.rx_in0
    .rx_in1           (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //           .rx_in1
    .rx_in2           (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //           .rx_in2
    .rx_in3           (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //           .rx_in3
    .tx_out0          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //           .tx_out0
    .tx_out1          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //           .tx_out1
    .tx_out2          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //           .tx_out2
    .tx_out3          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //           .tx_out3
    .test_in          (dut_pcie_tb_hip_ctrl_test_in),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //   hip_ctrl.test_in
    .simu_mode_pipe   (dut_pcie_tb_hip_ctrl_simu_mode_pipe),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //           .simu_mode_pipe
    .eidleinfersel4   (3'b000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          // (terminated)
    .eidleinfersel5   (3'b000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          // (terminated)
    .eidleinfersel6   (3'b000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          // (terminated)
    .eidleinfersel7   (3'b000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          // (terminated)
    .powerdown4       (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           // (terminated)
    .powerdown5       (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           // (terminated)
    .powerdown6       (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           // (terminated)
    .powerdown7       (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           // (terminated)
    .rxpolarity4      (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            // (terminated)
    .rxpolarity5      (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            // (terminated)
    .rxpolarity6      (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            // (terminated)
    .rxpolarity7      (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            // (terminated)
    .txcompl4         (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            // (terminated)
    .txcompl5         (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            // (terminated)
    .txcompl6         (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            // (terminated)
    .txcompl7         (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            // (terminated)
    .txdata4          (8'b00000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     // (terminated)
    .txdata5          (8'b00000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     // (terminated)
    .txdata6          (8'b00000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     // (terminated)
    .txdata7          (8'b00000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     // (terminated)
    .txdatak4         (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            // (terminated)
    .txdatak5         (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            // (terminated)
    .txdatak6         (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            // (terminated)
    .txdatak7         (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            // (terminated)
    .txdetectrx4      (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            // (terminated)
    .txdetectrx5      (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            // (terminated)
    .txdetectrx6      (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            // (terminated)
    .txdetectrx7      (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            // (terminated)
    .txelecidle4      (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            // (terminated)
    .txelecidle5      (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            // (terminated)
    .txelecidle6      (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            // (terminated)
    .txelecidle7      (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            // (terminated)
    .txdeemph4        (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            // (terminated)
    .txdeemph5        (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            // (terminated)
    .txdeemph6        (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            // (terminated)
    .txdeemph7        (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            // (terminated)
    .txmargin4        (3'b000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          // (terminated)
    .txmargin5        (3'b000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          // (terminated)
    .txmargin6        (3'b000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          // (terminated)
    .txmargin7        (3'b000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          // (terminated)
    .txswing4         (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            // (terminated)
    .txswing5         (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            // (terminated)
    .txswing6         (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            // (terminated)
    .txswing7         (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            // (terminated)
    .phystatus4       (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                // (terminated)
    .phystatus5       (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                // (terminated)
    .phystatus6       (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                // (terminated)
    .phystatus7       (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                // (terminated)
    .rxdata4          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                // (terminated)
    .rxdata5          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                // (terminated)
    .rxdata6          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                // (terminated)
    .rxdata7          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                // (terminated)
    .rxdatak4         (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                // (terminated)
    .rxdatak5         (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                // (terminated)
    .rxdatak6         (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                // (terminated)
    .rxdatak7         (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                // (terminated)
    .rxelecidle4      (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                // (terminated)
    .rxelecidle5      (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                // (terminated)
    .rxelecidle6      (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                // (terminated)
    .rxelecidle7      (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                // (terminated)
    .rxstatus4        (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                // (terminated)
    .rxstatus5        (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                // (terminated)
    .rxstatus6        (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                // (terminated)
    .rxstatus7        (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                // (terminated)
    .rxvalid4         (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                // (terminated)
    .rxvalid5         (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                // (terminated)
    .rxvalid6         (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                // (terminated)
    .rxvalid7         (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                // (terminated)
    .rx_in4           (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                // (terminated)
    .rx_in5           (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                // (terminated)
    .rx_in6           (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                // (terminated)
    .rx_in7           (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                // (terminated)
    .tx_out4          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            // (terminated)
    .tx_out5          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            // (terminated)
    .tx_out6          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            // (terminated)
    .tx_out7          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            // (terminated)
    .tlbfm_in         (1001'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000), // (terminated)
    .tlbfm_out        ()                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 // (terminated)
  );

  // The actual PCIe Hard-IP
  pcie_sv pcie_sv_inst (
    // Physical PCIe connections
    .pcieRefClk_in                 (pcieRefClk),
    .pcieNPOR_in                   (pcieNPOR),
    .pciePERST_in                  (pciePERST),
    .pcieRX_in                     (4'b0000),
    .pcieTX_out                    (),

    // Application interface
    .pcieClk_out                   (pcieClk),
    .cfgBusDev_out                 (cfgBusDev),

    .rxData_out                    (rxData),
    .rxSOP_out                     (rxSOP),
    .rxEOP_out                     (rxEOP),
    .rxValid_out                   (rxValid),
    .rxReady_in                    (rxReady),

    .txData_in                     (txData),
    .txSOP_in                      (txSOP),
    .txEOP_in                      (txEOP),
    .txValid_in                    (txValid),
    .txReady_out                   (txReady),

    // Simulation interface
    .hip_ctrl_test_in          (dut_pcie_tb_hip_ctrl_test_in),          //   hip_ctrl.test_in
    .hip_ctrl_simu_mode_pipe   (dut_pcie_tb_hip_ctrl_simu_mode_pipe),   //           .simu_mode_pipe
    .hip_pipe_sim_pipe_pclk_in (dut_pcie_tb_hip_pipe_sim_pipe_pclk_in), //   hip_pipe.sim_pipe_pclk_in
    .hip_pipe_sim_pipe_rate    (pcie_sv_inst_hip_pipe_sim_pipe_rate),   //           .sim_pipe_rate
    .hip_pipe_sim_ltssmstate   (pcie_sv_inst_hip_pipe_sim_ltssmstate),  //           .sim_ltssmstate
    .hip_pipe_eidleinfersel0   (pcie_sv_inst_hip_pipe_eidleinfersel0),  //           .eidleinfersel0
    .hip_pipe_eidleinfersel1   (pcie_sv_inst_hip_pipe_eidleinfersel1),  //           .eidleinfersel1
    .hip_pipe_eidleinfersel2   (pcie_sv_inst_hip_pipe_eidleinfersel2),  //           .eidleinfersel2
    .hip_pipe_eidleinfersel3   (pcie_sv_inst_hip_pipe_eidleinfersel3),  //           .eidleinfersel3
    .hip_pipe_powerdown0       (pcie_sv_inst_hip_pipe_powerdown0),      //           .powerdown0
    .hip_pipe_powerdown1       (pcie_sv_inst_hip_pipe_powerdown1),      //           .powerdown1
    .hip_pipe_powerdown2       (pcie_sv_inst_hip_pipe_powerdown2),      //           .powerdown2
    .hip_pipe_powerdown3       (pcie_sv_inst_hip_pipe_powerdown3),      //           .powerdown3
    .hip_pipe_rxpolarity0      (pcie_sv_inst_hip_pipe_rxpolarity0),     //           .rxpolarity0
    .hip_pipe_rxpolarity1      (pcie_sv_inst_hip_pipe_rxpolarity1),     //           .rxpolarity1
    .hip_pipe_rxpolarity2      (pcie_sv_inst_hip_pipe_rxpolarity2),     //           .rxpolarity2
    .hip_pipe_rxpolarity3      (pcie_sv_inst_hip_pipe_rxpolarity3),     //           .rxpolarity3
    .hip_pipe_txcompl0         (pcie_sv_inst_hip_pipe_txcompl0),        //           .txcompl0
    .hip_pipe_txcompl1         (pcie_sv_inst_hip_pipe_txcompl1),        //           .txcompl1
    .hip_pipe_txcompl2         (pcie_sv_inst_hip_pipe_txcompl2),        //           .txcompl2
    .hip_pipe_txcompl3         (pcie_sv_inst_hip_pipe_txcompl3),        //           .txcompl3
    .hip_pipe_txdata0          (pcie_sv_inst_hip_pipe_txdata0),         //           .txdata0
    .hip_pipe_txdata1          (pcie_sv_inst_hip_pipe_txdata1),         //           .txdata1
    .hip_pipe_txdata2          (pcie_sv_inst_hip_pipe_txdata2),         //           .txdata2
    .hip_pipe_txdata3          (pcie_sv_inst_hip_pipe_txdata3),         //           .txdata3
    .hip_pipe_txdatak0         (pcie_sv_inst_hip_pipe_txdatak0),        //           .txdatak0
    .hip_pipe_txdatak1         (pcie_sv_inst_hip_pipe_txdatak1),        //           .txdatak1
    .hip_pipe_txdatak2         (pcie_sv_inst_hip_pipe_txdatak2),        //           .txdatak2
    .hip_pipe_txdatak3         (pcie_sv_inst_hip_pipe_txdatak3),        //           .txdatak3
    .hip_pipe_txdetectrx0      (pcie_sv_inst_hip_pipe_txdetectrx0),     //           .txdetectrx0
    .hip_pipe_txdetectrx1      (pcie_sv_inst_hip_pipe_txdetectrx1),     //           .txdetectrx1
    .hip_pipe_txdetectrx2      (pcie_sv_inst_hip_pipe_txdetectrx2),     //           .txdetectrx2
    .hip_pipe_txdetectrx3      (pcie_sv_inst_hip_pipe_txdetectrx3),     //           .txdetectrx3
    .hip_pipe_txelecidle0      (pcie_sv_inst_hip_pipe_txelecidle0),     //           .txelecidle0
    .hip_pipe_txelecidle1      (pcie_sv_inst_hip_pipe_txelecidle1),     //           .txelecidle1
    .hip_pipe_txelecidle2      (pcie_sv_inst_hip_pipe_txelecidle2),     //           .txelecidle2
    .hip_pipe_txelecidle3      (pcie_sv_inst_hip_pipe_txelecidle3),     //           .txelecidle3
    .hip_pipe_txdeemph0        (pcie_sv_inst_hip_pipe_txdeemph0),       //           .txdeemph0
    .hip_pipe_txdeemph1        (pcie_sv_inst_hip_pipe_txdeemph1),       //           .txdeemph1
    .hip_pipe_txdeemph2        (pcie_sv_inst_hip_pipe_txdeemph2),       //           .txdeemph2
    .hip_pipe_txdeemph3        (pcie_sv_inst_hip_pipe_txdeemph3),       //           .txdeemph3
    .hip_pipe_txmargin0        (pcie_sv_inst_hip_pipe_txmargin0),       //           .txmargin0
    .hip_pipe_txmargin1        (pcie_sv_inst_hip_pipe_txmargin1),       //           .txmargin1
    .hip_pipe_txmargin2        (pcie_sv_inst_hip_pipe_txmargin2),       //           .txmargin2
    .hip_pipe_txmargin3        (pcie_sv_inst_hip_pipe_txmargin3),       //           .txmargin3
    .hip_pipe_txswing0         (pcie_sv_inst_hip_pipe_txswing0),        //           .txswing0
    .hip_pipe_txswing1         (pcie_sv_inst_hip_pipe_txswing1),        //           .txswing1
    .hip_pipe_txswing2         (pcie_sv_inst_hip_pipe_txswing2),        //           .txswing2
    .hip_pipe_txswing3         (pcie_sv_inst_hip_pipe_txswing3),        //           .txswing3
    .hip_pipe_phystatus0       (dut_pcie_tb_hip_pipe_phystatus0),       //           .phystatus0
    .hip_pipe_phystatus1       (dut_pcie_tb_hip_pipe_phystatus1),       //           .phystatus1
    .hip_pipe_phystatus2       (dut_pcie_tb_hip_pipe_phystatus2),       //           .phystatus2
    .hip_pipe_phystatus3       (dut_pcie_tb_hip_pipe_phystatus3),       //           .phystatus3
    .hip_pipe_rxdata0          (dut_pcie_tb_hip_pipe_rxdata0),          //           .rxdata0
    .hip_pipe_rxdata1          (dut_pcie_tb_hip_pipe_rxdata1),          //           .rxdata1
    .hip_pipe_rxdata2          (dut_pcie_tb_hip_pipe_rxdata2),          //           .rxdata2
    .hip_pipe_rxdata3          (dut_pcie_tb_hip_pipe_rxdata3),          //           .rxdata3
    .hip_pipe_rxdatak0         (dut_pcie_tb_hip_pipe_rxdatak0),         //           .rxdatak0
    .hip_pipe_rxdatak1         (dut_pcie_tb_hip_pipe_rxdatak1),         //           .rxdatak1
    .hip_pipe_rxdatak2         (dut_pcie_tb_hip_pipe_rxdatak2),         //           .rxdatak2
    .hip_pipe_rxdatak3         (dut_pcie_tb_hip_pipe_rxdatak3),         //           .rxdatak3
    .hip_pipe_rxelecidle0      (dut_pcie_tb_hip_pipe_rxelecidle0),      //           .rxelecidle0
    .hip_pipe_rxelecidle1      (dut_pcie_tb_hip_pipe_rxelecidle1),      //           .rxelecidle1
    .hip_pipe_rxelecidle2      (dut_pcie_tb_hip_pipe_rxelecidle2),      //           .rxelecidle2
    .hip_pipe_rxelecidle3      (dut_pcie_tb_hip_pipe_rxelecidle3),      //           .rxelecidle3
    .hip_pipe_rxstatus0        (dut_pcie_tb_hip_pipe_rxstatus0),        //           .rxstatus0
    .hip_pipe_rxstatus1        (dut_pcie_tb_hip_pipe_rxstatus1),        //           .rxstatus1
    .hip_pipe_rxstatus2        (dut_pcie_tb_hip_pipe_rxstatus2),        //           .rxstatus2
    .hip_pipe_rxstatus3        (dut_pcie_tb_hip_pipe_rxstatus3),        //           .rxstatus3
    .hip_pipe_rxvalid0         (dut_pcie_tb_hip_pipe_rxvalid0),         //           .rxvalid0
    .hip_pipe_rxvalid1         (dut_pcie_tb_hip_pipe_rxvalid1),         //           .rxvalid1
    .hip_pipe_rxvalid2         (dut_pcie_tb_hip_pipe_rxvalid2),         //           .rxvalid2
    .hip_pipe_rxvalid3         (dut_pcie_tb_hip_pipe_rxvalid3)          //           .rxvalid3
  );

endmodule
