--
-- Copyright (C) 2014, 2017 Chris McClelland
--
-- Permission is hereby granted, free of charge, to any person obtaining a copy of this software
-- and associated documentation files (the "Software"), to deal in the Software without
-- restriction, including without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to permit persons to whom the
-- Software is furnished to do so, subject to the following conditions:
--
-- The above copyright  notice and this permission notice  shall be included in all copies or
-- substantial portions of the Software.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR IMPLIED, INCLUDING
-- BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND
-- NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM,
-- DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
-- OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE SOFTWARE.
--
library ieee;
use ieee.std_logic_1164.ALL;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.ALL;

library makestuff;

entity rng_impl_tb IS
end entity;

architecture behavioural of rng_impl_tb is
	constant N                : natural := 1024;
	constant R                : natural := 32;
	subtype OutputType        is std_logic_vector(R-1 downto 0);
	subtype StateType         is std_logic_vector(N-1 downto 0);
	type ExpectedArrayType    is array(0 to 2*N-1) of OutputType;
	constant expectedArray    : ExpectedArrayType := (
		"11010010111000001100001110011010",
		"11111000100011011010111001001010",
		"10100100100000101110111001010100",
		"01010000010110010001010111011001",
		"01001100100001111101010011100100",
		"11011011100000000000100011101110",
		"00000011000011011010111100111001",
		"00001100100011111001011000001111",
		"10110000101010001110111011110011",
		"00100000010011100010110100100001",
		"10110011000010100000011000011110",
		"01101000010000011001100001101000",
		"10001001011000001110001101111010",
		"00001010011001101110110000010001",
		"01110100000110110011101100111101",
		"00000110010110000011001011001000",
		"11100110011101100011111000101101",
		"10000001110100101110001000000010",
		"00111011000000100111101111101100",
		"10001010011011011101000000011000",
		"00100001100010000101010101111101",
		"11001101010110000110010111110010",
		"01110000111000100110101100110110",
		"11010010101110111110101110000110",
		"01000011000000101000111011111001",
		"11111100110100011000101000010000",
		"00011110101101100010000110111101",
		"11010110000111101111110100100011",
		"01111000001010111010011010000001",
		"10100111110101111001000011000111",
		"11010101001000010011101110110000",
		"00001000011100111100000110011000",
		"10101010000111011111101000110000",
		"11010001111001000011101000000100",
		"11001000110000110101010100100000",
		"01101000000100010111001000110101",
		"00100100011000100111100001110010",
		"10000111000010000111011001011100",
		"10001010001110111011111000010000",
		"00011010101110000101011011010111",
		"01110000110001111100001001000110",
		"11111011100010000001100110010100",
		"10110011011011010011101000100111",
		"11111000101101001100001000111010",
		"00001001001001100000011100110011",
		"10100010110100100101000111010100",
		"11001011001101110000011011111011",
		"10110110010110100110000110111000",
		"11001100101110101110011010111111",
		"10100011011110000000100110010011",
		"01100000101100111010000111001100",
		"01010000100111100000101011100000",
		"00010111110011111000111010001000",
		"01011111001110101110100000011101",
		"01100001010001100010111110111101",
		"10010110111101001100000000101011",
		"11001101110101001111100110100100",
		"10100101001100001100101001011110",
		"11011111000101001010000101010110",
		"10010000100111100111111100011100",
		"00011111001100000000000101111010",
		"10010001111100101110010000100101",
		"01101110111011000010111111111001",
		"11100111000010111000010000101011",
		"00110000000001010010101010100001",
		"11111001111000000111000111011111",
		"10000010010000001010100011000011",
		"10010001010110110001110000101001",
		"00110000101001001001100111100111",
		"10010011110001100111011011011011",
		"11000011101101110100101111000011",
		"00001111100101000001111100010101",
		"11101110110110110110001001001101",
		"01100011110000111010110001100111",
		"10011100001001111000100011100101",
		"00100110110100100001111010010100",
		"10100100111001011111000111001011",
		"10001000111010001011001001101111",
		"00110011001011011101100001100110",
		"00011010101110100011010111110001",
		"01111100110011000000100100010001",
		"10101011001001110011000111101000",
		"10001110110100010011000010010001",
		"00111100001000010111111100110110",
		"11110001110110101000110001001010",
		"01110110000001111000011001100010",
		"01001111100011111010111101100010",
		"01100110001101001110111101101110",
		"11010110111010110100010011001011",
		"11101100110110111000101001010011",
		"11111111001001010111110001001100",
		"10001010001001110000010010110111",
		"11001001011101101011111011010000",
		"10111010001101011000100101100000",
		"11101110101011000010011000000011",
		"10000101101111011010110100001010",
		"11011111111111001110000000010100",
		"00011001010110000101000001011101",
		"00011101010010100110011111100010",
		"10011011010011001111011111101101",
		"01110011000000001001111101000011",
		"00001111110011001101111000001100",
		"00101010111101110011001011111000",
		"00100110100001100011011110010000",
		"01001001010100001000111011100111",
		"00000110100011110110111100000011",
		"10100100000011000010010010110001",
		"01001011010000001010111100111001",
		"10100010011110111101010011010010",
		"01011111011100101100110110110001",
		"00011000011110110001000001011000",
		"11111001110101110011011111101011",
		"00010110101011101100011001010011",
		"11110010101001011011001101010011",
		"11101100110010100101010111111001",
		"11010011110111110111111110001000",
		"11101011011011000010000010001011",
		"11110011000101100100001011001010",
		"00100000000100010011100001011110",
		"01000011101101000011100101010010",
		"00001001111010011010101001111000",
		"10001001000011001010011110000001",
		"01010100001001011010000111111011",
		"11100000010101010011011100100001",
		"01011001011101001100010000001010",
		"11110110101010011100110000101111",
		"10101110110001000000011101100100",
		"10001010011110100110100010110101",
		"10010001010110001110001111001010",
		"00000100101011010011000111101010",
		"01001000011101000011001100100100",
		"00010000001101111101000000000100",
		"10010101101110011101000000000100",
		"00010001001101111111101101000001",
		"00011000001010110001000111000010",
		"11111001011010010111010011001101",
		"11011001111110000101010101110010",
		"10110000110000110011101000011100",
		"11100011000011010001110111000111",
		"01001110110001111100011100110000",
		"00000010010011110010010110001011",
		"11000110000110100101110010111110",
		"01001001000111011001000000001010",
		"00001001100000010010000001111011",
		"11101111011010100101101101011000",
		"10101110100110111000100001101000",
		"10010010100110101110010001010100",
		"01000110001011101101101001011110",
		"01011011100110010001011110001110",
		"00010110110011011011111010111101",
		"01001110011110101010010000111111",
		"00011100101110011011101010011101",
		"00000101111011110000010000110110",
		"11011111111110001110101011011100",
		"11111000111001010110000110000111",
		"10110100111100111010001100001100",
		"11101111001110101111111110001110",
		"11001100000001000110001111010110",
		"10000111011111001111110100101101",
		"11111111000010010111001101001101",
		"00101101001110001010101101000011",
		"01011111000000000110010110001100",
		"11100011111111000101011011100101",
		"00010001000100111101000111111010",
		"00101001010011001110110110000101",
		"11010000111110110111100000100011",
		"11111010011000111000101011101000",
		"11100010010110100101001101011101",
		"01101010100110001001110100010000",
		"10110111111000111001011101100010",
		"11000111001001111000010101001011",
		"11011101100011010101001110010001",
		"00111010010101011010110010001110",
		"01101111001000111010000100010111",
		"11111010100001011111010000000110",
		"01111000111000101100001100011100",
		"00011010100001001001101110111110",
		"00100010000110001111110000111111",
		"11111010101000100010100001000010",
		"10001110101101000011000111110100",
		"11100000011001011100000111110101",
		"10010010110010101111011001000110",
		"10101011100001100010011111001001",
		"00000101101010010000000100101010",
		"11000101000010010011101001100010",
		"10010011101011000110100110000000",
		"00011011001101101110101100101001",
		"10001001100101011011110000000101",
		"11010011010100010101011110110001",
		"11000111010010110110100101010001",
		"11110000001010000101011111110110",
		"00010100101111011110001111000101",
		"11010010010100010011101101110000",
		"01100011011111111110011101000011",
		"00010111111010101111111000001001",
		"01000011101110011111100101011000",
		"00101111101110101000011010100001",
		"10011000100110001100110101001000",
		"11000010100110010001011100001110",
		"01100010110001000000110010111000",
		"10110111011001000111001001110110",
		"01001000000001100111110001110000",
		"00011000111101101001010011001001",
		"10101101111111000010101010100010",
		"11101111010100001111110010011101",
		"00100011001110111111101110101001",
		"11111010001111111010010101100011",
		"11110011001011011000111111111010",
		"00101110001010001100100010100001",
		"11001101010001001101011100101010",
		"10011111011001010010000000110101",
		"00011110010011010111011000101100",
		"11110100010101000010100001001101",
		"11101001111010111011101000111110",
		"11101011001001111101110011110000",
		"11000110111110100001010111100011",
		"01100100110001011001100100000010",
		"00100010010100011010010010100011",
		"00011110111110111000110001001011",
		"00001111010101110110000111111110",
		"10011010110101000101001000010110",
		"10011001100110000010010000111000",
		"10111111110010101001011001110110",
		"10000001001000101101101001101001",
		"00011110001011001010110100100011",
		"00100001011010010011111001100100",
		"11000011100111001001100001011011",
		"11001001001001111011011111010011",
		"00001101000011011110000111000100",
		"01010111000111011001100110110110",
		"10010001111000101010011001000101",
		"00000000101010101001110001100011",
		"01110110111001011110101111101000",
		"11110100110010010000010000100111",
		"11111100000000010101110110011111",
		"10111001100011101000011010100110",
		"11010100100001000010011111010110",
		"01110101111100010011100110010000",
		"10000110010011001110111000110000",
		"10110110011101011001000111100101",
		"00111110111110100100111101010110",
		"11011101010010001010000001101010",
		"10010110001010101100100001000001",
		"00001000111011101100110000011110",
		"11010010111101100110101111000101",
		"00101000111010101011001101100111",
		"10000100110110110000001000000010",
		"11011001000111100111111111111111",
		"01001101101011000001111100110110",
		"11010110101010011101000101110001",
		"10000010100101010001011011111001",
		"00011110001110000010001000011010",
		"01110000110100001010111001111010",
		"00101101010110001000000010001101",
		"00001101011010010011101000001101",
		"10101100000011111011100011000000",
		"10101010000111101011100111111100",
		"01111100001111001110100111010100",
		"00010101000001111001011100111100",
		"00101010110100011101110111000000",
		"10110110100000011101011111111011",
		"00100101101010011101011100101100",
		"00110110110110000101000111010000",
		"11110111001001000001000111101111",
		"01010100011110011101100100010110",
		"10101101101111110111110011000001",
		"01001110110000000110101110111110",
		"01101110000011110010100010111111",
		"10001010001101000010010000100101",
		"00000001010111001110010001101100",
		"11111010011011111101110110011111",
		"01011111110000011000110101010010",
		"11000000000101010000110101110010",
		"01001010111101000011101011111001",
		"00110001110001111100010111001010",
		"01001000000110010101110011010101",
		"10111010000111110100101010101111",
		"11101110001110001111100010101110",
		"11111010010111100101011101111001",
		"00001011010011010010010001010101",
		"00010011101100001000100011011001",
		"01111111101111101111100111101100",
		"00011000010110101100000011101110",
		"10010111110000001101100110001101",
		"01010010111000010101100000010011",
		"11101101110110011000000101000000",
		"00011001011000010001110001100011",
		"10000010011000011000001100001111",
		"10101010010110110010000001011110",
		"00011010111100001100100010001000",
		"01000100101100011101001111110111",
		"01010111011111010011011010011010",
		"00001000100010001001110111110011",
		"11010010100001010010100010101110",
		"00000000100100110100001101110110",
		"10001010100001101011011111011000",
		"11111111110010001111010000101001",
		"01110100010011101001101100011110",
		"11100110111001100101101101001111",
		"00100001000010010111111010001110",
		"10010110111000000111010010001011",
		"00110100001011100111100101010000",
		"01101100101001011101101010101100",
		"00110101101101111011100011011001",
		"01111110101011100011011101010011",
		"00110000000010000101001011101000",
		"00010100011010010110010011010110",
		"00100010011101111001010100101000",
		"10110011010100110101011111110011",
		"11101110110010000010111001100000",
		"01001110011100010100010110000101",
		"10111111111010010100101000001110",
		"01010011011010010001010011001011",
		"00100100101100001011100111110110",
		"00000001110110010011001011100100",
		"01101110010101101110101110000011",
		"01010010001000111000001001110111",
		"11101111001001011000000001100000",
		"10011111101111010000110110100111",
		"00101110111001110001011011111110",
		"00000010101001000110111011100011",
		"00011001010000000000000010110000",
		"01001111001100011110011111010100",
		"01110001000100011000111100000000",
		"10100111110100000111100001001100",
		"01101011111001111000011111011001",
		"10100000100111100111110010111110",
		"00011111001011010111100011000011",
		"10011100000101110101111110101000",
		"01010011101100111011110111100000",
		"11110010111001010101101110000101",
		"10100000010110011101001000011010",
		"11110111100101111010111101111010",
		"01001100110111101000100101101110",
		"01000100100001000001100010101110",
		"10001100001000111001111110011000",
		"00000100110001100110000001001001",
		"10101000110111010111000110000101",
		"00111101101010001100100100110100",
		"10110010011011011101110011100111",
		"01000000000101100111000101101110",
		"11000110100110111001110011100110",
		"01010011010001001011100011101110",
		"11100010101010000101100100101100",
		"01011010010010011110111100101111",
		"11111101010010010100111110101010",
		"01100011000100011101111100011110",
		"01100110100010101111010001111001",
		"10010010101000100000111100111101",
		"01101111110010001010100001111110",
		"10110110101011100110100000100000",
		"01100010001111010010111101111110",
		"11110100110101100111001001111110",
		"00000100100001000000001001000010",
		"11111000101101010100110111100110",
		"00100111111000001101101101010001",
		"00010001101111110011101100010100",
		"11000101010001001100010110101011",
		"00001101010011101011010000111000",
		"01101100100100111010110001000011",
		"10001110100100100111111100111101",
		"11100000010101010001110001000111",
		"00100111010101001111100100100100",
		"00011000101000000101011011010011",
		"10001001011010101010000110010111",
		"10111001100111000001001111110110",
		"10001001001100010010011001010001",
		"11011110010000001001001011100001",
		"01000101010110011000000101001110",
		"00101001001101111101010111011011",
		"10000001011010011111110000110100",
		"00010001111101000010011010010111",
		"00111000110100110000010101011100",
		"00111100010001101001000000100110",
		"01100000010001111000000100000010",
		"10100100000010100110010110011010",
		"11110100100111011001000001011001",
		"01001001101001111010001011111001",
		"00110110001101010111111011110110",
		"01110101111101011000011101011100",
		"11000011100110101101100101110011",
		"11010011111000111011100010100101",
		"01010111101011010110001100000001",
		"00000100010011001111001111111111",
		"11110011100000101111111100110011",
		"10001011010110001001000101110000",
		"00010100000011111010010110010100",
		"01001101011100010110101010010110",
		"01100001101010000010111100000101",
		"00101000010000000101100111101111",
		"01100111111000101100010011111001",
		"00111101001000011001111100110100",
		"11000001101010101111010011000011",
		"00110010011000101110110011000111",
		"01111100001011110011010110110001",
		"10101011110000000111011100011001",
		"10101010000100100101001100011000",
		"11111111101110100101100000010001",
		"10000101000101101011100101101101",
		"01101011111001010111110110011000",
		"11000001101011101000011110111100",
		"00110000011010011000011001000101",
		"00011000100100110000111000110001",
		"10000101001100100000111001100010",
		"01111000110001110100000111010011",
		"10001110101101011011101110000111",
		"01101000101000111001100100100000",
		"11001011001101000101011101100011",
		"01101001100101000010110101011010",
		"00100101011001011101111101011101",
		"10101110111001101101101001111010",
		"00010001001010000000101111111110",
		"11111010111010000111010100000110",
		"10101100001011010100101100101011",
		"10001110011001111100100110000110",
		"01110011010110100110111010110010",
		"10111101001010001100010101000100",
		"11111000000111100011100110000010",
		"11100100101110110110001000100110",
		"01000111100011011100111000001110",
		"00011000000001100101000111111000",
		"11110100000001010001101000010101",
		"00010110111011101101100010100100",
		"01010100101111010000111101101001",
		"10000001001100110000101000111011",
		"11100100000110010110100010000100",
		"11010100101101001110010110101110",
		"00011111110100011101010110111000",
		"10100000110000100000100101010111",
		"00010111010011110110101010101111",
		"11011100101010011010111011101010",
		"10111101000111000010011101100011",
		"11010110011100100000101111101101",
		"00111001111010101001111011001011",
		"11101001011010101101010100000111",
		"10111001000100011001011101110001",
		"10001001111001110110011011100111",
		"00010010111110000000110011000111",
		"10101010001010111110000100110101",
		"10011101111101100010101000010001",
		"01101010011111110011010111110000",
		"10010110010111111000101100000111",
		"00100001001010001010111010001001",
		"10011101101101110100100001110111",
		"00110000100000010100000011111111",
		"11100110010000000010010111110011",
		"01111101100000011101000111101110",
		"11101101111111101001111001011010",
		"00111101110001101101010001101001",
		"11111000010100000100001110010100",
		"01010000001011100000100001000110",
		"00111100011011010101011101110011",
		"00011110110000001010010111010000",
		"10011000110111011101000100000100",
		"11000111111011001001111111010110",
		"10000100110010010100101010001001",
		"10101100001001101001100011111011",
		"01011011000001000000010011101010",
		"00111000010011100011111111011010",
		"11111011001010111110011010111011",
		"11011101100001101101110011100010",
		"01001000001110000110110001001000",
		"00100110001001000001001100000000",
		"01001111111010111001111100010101",
		"11010001011101101011110010001010",
		"00000111110000101111110000000110",
		"01010100011100111100100101000111",
		"11001110011100100001111100000001",
		"11010110110110110010010001010010",
		"11100100001100100011000010101100",
		"10100101111000101001011010110011",
		"11010011011000101001111001001000",
		"01010000101000011101110111000111",
		"11000001110100101000000111001001",
		"10111110011011010110111100001100",
		"11001001001010000000000110100111",
		"00101100111000100011011010110111",
		"11111100010000001110001101110010",
		"10110010010100111010000101100001",
		"11001110111011101000011001110111",
		"11110011000101110101001110110100",
		"00101011011100101010011011010010",
		"10110011000111101100110011011101",
		"10011010101111000010000011000000",
		"01010000011001110000010010000100",
		"00110101111101001100010000111111",
		"10001110110111001010110001010010",
		"00000100011111010000101101011000",
		"01010100010101000100111001000001",
		"00001001000101000101110110010111",
		"00000001011110100001011001001001",
		"01111011000011001011011110101110",
		"11000010100010001000010001100101",
		"00110100111101110001110110011001",
		"01110110010011001000110100100000",
		"11010010101110000010001110010100",
		"00000111111111100100000111110001",
		"10011010010000010000100001000000",
		"10101101101000000011001000100011",
		"10101010000000001110110110011011",
		"10010001001000001010110110001001",
		"10101111101101111000111010111111",
		"11011110101101110111001000001001",
		"11010110001000111011110001010010",
		"10101000111100001011110111111010",
		"01000011110010011111010000000110",
		"11100000000100011100001010111011",
		"11011111101111011000110101000101",
		"01010110101011111110011111001101",
		"01111100001111101101011011010001",
		"11011110001011010000001100101001",
		"11011101010101000011101100000101",
		"01110110010110111110100110100110",
		"11001110100101010101011110010000",
		"10010111101000010100110011011000",
		"11011011101011100001010100010000",
		"10111110011010001000101001000010",
		"00001010011011010011111100101111",
		"10001010001011000101101011110000",
		"10000111011110110000101011110101",
		"10010101111110100100101111011111",
		"11010000011110010000110100011010",
		"11110100000100000101111011010110",
		"00110110011100010011010010001000",
		"10000000000000110100111001111001",
		"00101001110001000110101001001010",
		"00000011100101000110001110000001",
		"10101010001100111101110110100011",
		"00101101010111110011111011000000",
		"11110001011011110101101101010010",
		"10100010000010100011001111100111",
		"11111101010011101010011001011111",
		"01001011110010010110011101100111",
		"01100101110100010100010000000111",
		"01000111011110100111101010100110",
		"01011111010100000101000101000101",
		"00111111110010011010010100011011",
		"00110000000111100000100110110110",
		"11110101100111110111110101001110",
		"00001111000010000001111010011001",
		"00101011101000101010001111110100",
		"01110001111101001110000011011100",
		"01101011110111111111100011110011",
		"11000011000010001011100011111011",
		"00000000111000110101110111110010",
		"01000110100011011001111110100010",
		"01011001010100001111111010110001",
		"00001010111001011110011010100010",
		"10001010001011111111101010110010",
		"11000011101100111001011000010011",
		"10110101010100100000101110110101",
		"11100001101000001101000110010111",
		"00000000001000000001000100001010",
		"10000101001011011000101011000111",
		"00011011010010010010010101010111",
		"10000000010010110010111000101101",
		"11110100110101010100110000101011",
		"11001101110000101111110111001011",
		"00111010010010001010111101111111",
		"11110110111110001111100000110000",
		"11011001011011111001110111000011",
		"11001000111011101111001000011011",
		"11110010101011110010100000000001",
		"00000000110000001100010001111111",
		"00001001110001101010110101110111",
		"00010011111011000101110100100010",
		"00010011011011110011000010001001",
		"00000101001100101101011100001011",
		"11000110111111001111011010100110",
		"01111010001000111001010010001011",
		"10100100001010101001101000100000",
		"10011011011101001100111011101100",
		"00110001100100111110000011111111",
		"10000101101000000101100011000001",
		"10000001101110100101001001011011",
		"01100101110111111100001001100000",
		"11010111111001010111010101101100",
		"00001000001011010101011001110001",
		"00011101101100010111001110000100",
		"01101111111001000011101111000100",
		"10000111101011001001011100001111",
		"11100000100100100000010100000000",
		"10101110000110011101011100011111",
		"01100001110101101000000111111011",
		"00000111111001010001111100110001",
		"00001011000101101101101001011001",
		"01011101000010010101011001010001",
		"10011100100100011000100000010010",
		"11001110100101011010011100100101",
		"11010011001000000110110101100011",
		"10100000111011101000111010010000",
		"01111101001010101000000101101001",
		"10111101100011001111111100000000",
		"11111000010001110001111011010010",
		"11000011010101111100001010011110",
		"00000110101111011100111111110111",
		"10110001100000000100110100111001",
		"00011101000100000000111000001011",
		"01111001011001000001110100101101",
		"00110101000010110101110011000101",
		"10111011110110101101011100110111",
		"01110110111011110110100100000011",
		"00101001111001100000101100100100",
		"00011110101011100110100011101000",
		"01001010010111011100101010101011",
		"00011000000011001111011101110011",
		"00111111001000000000011101001100",
		"11001101001000100011100101000010",
		"00101101000110101001010100000011",
		"11000011000110100110101111001000",
		"00000000001111100111001010111110",
		"11111010100000100110100111001110",
		"00101010011111000011010001001110",
		"11100111011100110011001100010011",
		"11000110110011111101110011111101",
		"00100110110010100000010111001100",
		"10000111101111101111001101101010",
		"10010100100110010111001101000001",
		"10111110011100000010000101001110",
		"11111010100110101010000101000000",
		"11101110100110110000111010111101",
		"01111100001001001100101000100101",
		"01110111000101101010010011000110",
		"00011010011111110110111010110101",
		"00001010101101100001001110001001",
		"11101011100111000101001000100001",
		"11010110000010110110101001011000",
		"11101001100100111101111001011001",
		"10010100000010011101011001101010",
		"01110000001001001000011000111001",
		"11000011111000001111110001001101",
		"01111100010011001001101100111111",
		"01100001010010101010110101110111",
		"11101100011010010001010011001011",
		"10000011110111011111011111101110",
		"00111110100010111100110001110100",
		"00100010101011101001101011100010",
		"00011010001001001010010001011111",
		"10100111001001110111011110111001",
		"11010101111011110010001110110100",
		"00000000111100011110111010110100",
		"11101011011001111101100011011101",
		"01110101011100011010010011111001",
		"01100101010100101011001011001111",
		"00010011011001011001101001001010",
		"01111100100100000010111101011110",
		"00110111110010100100101110111101",
		"01001110011001101010100010001010",
		"10110001010111010100101001010000",
		"00111001111000111000011101001000",
		"10001010110010000100010101110110",
		"11011100001001001101000101101011",
		"00011110001011111100010011001001",
		"11110110111111100101101010001110",
		"01110001000010011101000001100001",
		"11011011011100001000110001010001",
		"10010000110011001101011011110000",
		"00100011111000101100111000010000",
		"10010010110111000111010100111100",
		"11011101110101111010111000100011",
		"00100001100111111110010011111111",
		"00100001101110111000000010001111",
		"10100000101010100101111011010001",
		"10101101000001001011010001011110",
		"11111000010010000100011100111110",
		"00000010001100100100001001110001",
		"01011000111111110011011100000001",
		"01000010111111101001110001000001",
		"01010100111011000101100100110000",
		"00100110010100110001010010011110",
		"01101010011100111111101110010000",
		"11101010010010100011101001100110",
		"01101000101001000100110000001100",
		"11110011000101011110100011100101",
		"01101011011001000100111000111101",
		"00100001110101100100011101100100",
		"11111011001001011100101110000110",
		"01110000101001110011111011001011",
		"10110000111100110011101110100010",
		"10100100110000001101010101110100",
		"01001000111000110111001010110000",
		"11000101010101100101111001100100",
		"01111101000011010101010001110010",
		"10010101010100010000110000101110",
		"00011010010110110010110100111101",
		"00010000111000111011011011001110",
		"11000000000010000010110101111011",
		"11001000001101111111010010010101",
		"01001101110000100101110101110110",
		"00111011110001100010011100111111",
		"01011000000010110111010010000111",
		"01101101000110001101100100010110",
		"00000001000000100100000110011111",
		"10110010110110101111100000000100",
		"11001001011001100111001011100110",
		"00101101001111111001011110110100",
		"11000010010100001100110011011000",
		"01000111010010001010101010001101",
		"00000010100010111001011111110100",
		"10000011010001011101000111110000",
		"01001010001111001001110110111010",
		"00000001010011011001000011000011",
		"10101111111111111000111101110001",
		"01001111100111001101101111111010",
		"00110101011000100001100000101110",
		"10000100000110100000111000000100",
		"00011010110111100000111100110101",
		"00001011101100001011011011100010",
		"11111011001000101110011110101100",
		"00000101111110100010001100001001",
		"11011111010110001000110001000011",
		"00111110011010011011000010100111",
		"00010110100001100011110101110000",
		"10000000110111000000010101001011",
		"00111101110100000010110010000001",
		"01000010010110011101000111110100",
		"00110111010101000111111100011101",
		"10010010000000011110001001101001",
		"01011000001101000000001001011100",
		"11111101100001010100101100010010",
		"10111001011010011100110001011110",
		"00011001010011010101111010111110",
		"01101110000110001100011110001100",
		"01101110011001000110011101111011",
		"01101000000011100100010110100011",
		"11001110100010100101100110100100",
		"10010111111100011111101001100100",
		"01111001010010100011001111100100",
		"01010111110010010110001110100011",
		"10011100110011010111101100110000",
		"11001111000010101001011000111001",
		"11011101000010101110011100010011",
		"00110001111100001010110101000001",
		"01000111110001101001010110001110",
		"10100111001010010100010110100100",
		"11000010100111111101011111010101",
		"10110011010101101110010101010001",
		"10101010000011011001100010100001",
		"11101001011010101001001010101011",
		"10001101000000100101101110010010",
		"00000110010110011010011100010000",
		"10001111001010100100111000000101",
		"11001111010101111100000010000001",
		"11000100000000111101000110011011",
		"11110001110011110010110010101111",
		"00011011010100001010110111000011",
		"00110010111111000100001000010110",
		"00100011111001010001011101111101",
		"11110110110110111010101011101001",
		"01011110100101100001111100110110",
		"01000101111011000000001101101011",
		"11000001101110101101101110010011",
		"10110100000111001010101000111111",
		"11101100100001111011010100110011",
		"01100011110111100101111101110000",
		"11010000100001001101000001111000",
		"11111100011100010100101000000000",
		"10100011111000111000011001110111",
		"01010001011111100010100010101110",
		"00000100010011100100011010011010",
		"01010010110101001011011000011000",
		"01110001100110010000101101010110",
		"01100110101111011110100111010101",
		"11111000110000101101101011010110",
		"01110011010010110101101000010111",
		"01111101101010110010010100001011",
		"10010011011100001111100101011010",
		"00100010000101100011011101001110",
		"11001010100110110010011000001110",
		"01001111001100001101000101110010",
		"01000011011101001101010111000111",
		"00101101010000111001011110011010",
		"00100110110010000111100001110000",
		"00111101001011110111000101101100",
		"01000101110110010011110011011010",
		"11110110101001100001001000011101",
		"01110011100001111110001010111100",
		"01011110010011101010110110001011",
		"01101001111110101001100101111101",
		"01100101010001101100100110101001",
		"00000000100111101011101000000011",
		"00001110110100110001000101111110",
		"01101000010100111000010010000000",
		"10011010010001001010111110011110",
		"00010010111100110100010000000001",
		"10010110101111100100110001110010",
		"01001101100001000011010001010000",
		"01110101001100111111110001111110",
		"00001100100001100100000110010111",
		"01001110101011001110101101101110",
		"00011000100100011100001111010001",
		"10011110010001110000100101001110",
		"01110111011101110010011111111111",
		"11011110010110010010110010000000",
		"00001010010001110101010000001001",
		"10100111001001111001110110010001",
		"11000110110110110000010001010111",
		"11111101010100110100011001010000",
		"00000010101101000011010010000100",
		"01100101000001000011110100011010",
		"10100110111010001100011001100100",
		"10111010110100001000110000101000",
		"01010111100100110110100000101111",
		"10110111010100110110101000011000",
		"11001001010001100100001111001111",
		"00100000000000000110100001101110",
		"01110101000010111011100101111001",
		"01001010111110100000010001111010",
		"11110111101010001011101010001000",
		"01011010101010001110001010001000",
		"11000100001001101111111111001110",
		"10110000101100111110111010001011",
		"01111010111111001011011111000000",
		"10111110000011000001010111111010",
		"10010111001011010101111010111100",
		"01110011101100010011001110100110",
		"01011011001011001100110011010000",
		"10100110001001111011001011111110",
		"10001101010011100011011101011110",
		"01100101001100000001111100000101",
		"01100110101010000111001111101010",
		"01110110110010010010110111100110",
		"11011001110110101011110000111100",
		"00110100110010101010000010000111",
		"11011100010000001111110010011110",
		"10001001100101011000001111001000",
		"00011101110101001111001010100011",
		"01000100101100010101111111010111",
		"01101100110101010011010011011000",
		"00100110000001101011000001010101",
		"11000100010110010011010000111110",
		"10101001000101111001101000010111",
		"10100101101010110111110110101110",
		"11000011101001010001110101100011",
		"11000011001111000110111101111000",
		"11101100000101101011000010100010",
		"11110110110111001000100001001011",
		"10110010111010101101001100101111",
		"00001110101100001101010110011011",
		"00110101010011110000011000000110",
		"11001101100010010110011101101011",
		"01011110100000100011110110010001",
		"01101101000001111100111111000010",
		"10111101000101110001000001110110",
		"01111100110011001010111100010100",
		"00011101010101111100110101110010",
		"00110100100101101010100011010001",
		"00000001100010101100000001011001",
		"10101101110000110000001111110011",
		"00011000111001010010101010010100",
		"01001100001000110100011110101111",
		"00100111000001001000110001011011",
		"00010110000111110101000010100000",
		"01100001110011111001100001100010",
		"00101001111001011110000010000001",
		"10101011100010010111001010101011",
		"01100110000010010111001110101000",
		"11001100000101010001100111010001",
		"00100111111111000010000110110110",
		"10101110100000101011010110001011",
		"01101010100011001110100101010000",
		"10001110101000101100111111101100",
		"01110010010111101110111000011010",
		"11001011011000110010111010100100",
		"10001010100000111100111110000001",
		"01101110110100000001100001111110",
		"01000010100001111101110111010001",
		"10001111100010000011101010111101",
		"10010101000110110010010100001011",
		"01111000111111000001010111001011",
		"10111011010000100010110011011011",
		"10101111101110011010111001011110",
		"01010000000100010010110000101111",
		"00101010000101010011010111011010",
		"00101010001000001011101100001001",
		"10001110100010000011000001110001",
		"11101100011011100001111011111110",
		"00100100111101001001010000100110",
		"01110010011000010010001101000100",
		"01111010001111000000111001111100",
		"10100010000000001101000001100100",
		"00010110011100010001101001010110",
		"11110100000110000111000000011101",
		"10111001011101100100110100011000",
		"10010110000010100010000001001010",
		"10011011100110011100000010000101",
		"11010011010010000100010001111101",
		"10010101110111001111011111101000",
		"10101111111100000110011001010000",
		"01100010111010011101110000100101",
		"10111100001011110100001100110110",
		"01000100111111010111111100001001",
		"01010110010101001110000101110101",
		"10101011111001100011111100101010",
		"01111001010111101101010001111010",
		"11011101001000010110110000010111",
		"10111100010101111010100110110001",
		"01000011010010010110110100100100",
		"01001111011101111000111110111101",
		"10100000011100010000111111001111",
		"00110001111000100111011000100111",
		"10001000100101000101010001101011",
		"00011011110001001111110100010101",
		"10011110001100101101100111110110",
		"00001101101011001000011110000110",
		"11010110000111011100110100011000",
		"11110011010011001101100001110000",
		"11011011101011100101010010101100",
		"10100101110010001101101001000111",
		"10001110101101101000111001010011",
		"01100111100001100111011001101001",
		"01001110100001000011101011000111",
		"11100111110100110011100011101101",
		"10111001100011111001010111010000",
		"01110100001000011011110101011010",
		"11001100111101011010011100010001",
		"00010100111011000110101001100000",
		"11100011001100010110110010110110",
		"01111100100111010110101001101100",
		"00010001001110101001110001110010",
		"01001011011101101100000001001100",
		"01111110010001101100011111010100",
		"01010001001110001101110000100111",
		"10001111110010101100010001011101",
		"00000011111110110111101010101001",
		"10010010010100011011000110101101",
		"10011001010111010000100100011111",
		"11001100010110110111100001000000",
		"01100001100110101000111001000011",
		"10110101101000111110111111101000",
		"00011100100010111010011001111110",
		"10001101100001110110011100110010",
		"11010011000100110000111110100100",
		"00011110111010101110010101000101",
		"00001000110010000001100101001001",
		"11101011010110011110101011100001",
		"01010101010000100100011100011111",
		"11001000101110100111010011111110",
		"11011001001100001011101110010100",
		"00100011010001001101000110110001",
		"01101110110111100010100001001111",
		"01010100101010010101110101111000",
		"01010011100000010111100000011100",
		"01010100101000010000010110010000",
		"00011011010110000000100000011111",
		"01000101010111011010011100000111",
		"00000100011101010000010100101110",
		"10001100111011101110011000100001",
		"01000110110111100110110010010111",
		"11011100110010100010101110011000",
		"11111010111011001111110010101100",
		"11011111011011011001010000000001",
		"00100011110010000100000101111101",
		"10110111100000000100101001111100",
		"00011110111110000101101000111100",
		"10110010101011000011010110101011",
		"01000010100011110101001000011110",
		"10011110001010100100110010000010",
		"01001100100011100010000001011001",
		"11000011001010001110101110001000",
		"10001010101011111101001110111101",
		"01100111101100010110111001101100",
		"10101111011001001011011010111100",
		"00000101010111101101110100010100",
		"00111001111110000000001011010011",
		"00111110011110010010101101000010",
		"11110110000001111100111110000100",
		"00001000001001110010100001001101",
		"00010110010001010011110111100111",
		"11001010100101111010001100001010",
		"11110000001000100001001010100111",
		"01001001000001100101100111011100",
		"10000101100000011011011100110111",
		"01101010000001010000101111111000",
		"01111011111010111100101110000101",
		"01010111011001001101101100011001",
		"00011100110110110100101011010100",
		"10010100111101010011010011111110",
		"01101110010011111011111101111011",
		"10010001000110100110110111110110",
		"01101100110010101000011110111011",
		"01011100110100111100001101110111",
		"00101000011000111110101110000011",
		"10000001111111111010101001011100",
		"10110111000101000101011111110110",
		"01111010100011001101110001101101",
		"01110000000010010001001101001101",
		"11000101011010110000000101101000",
		"10101101011111110101001011001010",
		"01101000000111000111101011101011",
		"01011000001000111000111000011001",
		"11010001101100011010010000000001",
		"11111000111010010001000011001001",
		"00111110101101011010000010100010",
		"01111100010000011000101011000101",
		"11110111100000001101101010001001",
		"11101100001111010001011001011110",
		"00111101010111001101010100000110",
		"10100011111111001100100111110110",
		"10101101111101000110110011010001",
		"01100011000100101010000011110101",
		"00110000000010101000001100000000",
		"11010111110010010111111001000110",
		"10100111100011111110001010001111",
		"11100000001111000001101001000001",
		"11001101100110010101001101011000",
		"10110110110101101011000000110010",
		"11011101110011100001110000010110",
		"01110111100101110110101011001000",
		"01111011110000101011001011111000",
		"00101010011111000011111001001000",
		"01101011111101100110111000100010",
		"01011011101111101001011110100010",
		"11001101100111010100001010000011",
		"00001101000010000000011001101110",
		"11101101101111000111010001010101",
		"01101011000101010110101010111110",
		"11111100111111111010000101100011",
		"00111000000110101001111101001010",
		"11001000100111110010101111110011",
		"10111111000001111101110100000110",
		"01001010101110110010011001100000",
		"11000010100001100010111001010000",
		"10010100110001100110101010111101",
		"11001110100010000101111111001001",
		"10010010001001011111111001001001",
		"11010011111001001111110000100000",
		"10011001011010001011101001001011",
		"10010110010000001101010101011100",
		"01101011011101111110111001001000",
		"10000001100010111011110101101101",
		"11011100011000011010101101011001",
		"00011011010001011111111101110100",
		"00101001100010100001000100101000",
		"10100111111100011100010100100000",
		"11000000000001101010110001000000",
		"01100010100100000101001011011001",
		"01100010100110100010001101110110",
		"00000000110010100010001000101001",
		"00000100101101011001010011110010",
		"10100111001011011111111001111001",
		"10111100111001010111001010001011",
		"10000101000110000110000100001101",
		"10001001000001101010111000001000",
		"01000110000100011010101011101010",
		"11101010001100000010000011000010",
		"00100010011111001001011100101101",
		"11001100000101100110000001100001",
		"11000100100001111110000101110011",
		"11001101111001101001000001000010",
		"01110111001111100001101101001110",
		"10001101111110011110100000010000",
		"10100110110010111000101011010101",
		"11011111100101101011011011110100",
		"11000000010010011000110000111000",
		"11100101011001100001110110011010",
		"01101100101000110010010101011010",
		"11111111100100010000101000000010",
		"00110000001001010111000110011011",
		"01000111010100100100111110100110",
		"11001010001000100111000010110011",
		"01101010000011111111010110111001",
		"11001110101111000111100011100111",
		"10101010011000101001101110001000",
		"00001001000100011111101001111111",
		"00101101000100001010100011100010",
		"00101110010011101111110001110111",
		"01001100010110011111011101011101",
		"01001011010001010100110000101110",
		"00101000011100010110101000110110",
		"10010011100011001011101011000101",
		"10111111110010001010100110011000",
		"10011001000010110100101010111010",
		"10001101001001101000000111000101",
		"10100101000010011101110010100101",
		"11001011011010100000110111100111",
		"11011111000000111111110011001101",
		"11100011001000111011101011100000",
		"01001001010101001010011100000011",
		"11101111101011001011101101110010",
		"01000100100010000111001010110111",
		"11111110100110010011110000110001",
		"00000111100110110011100011111111",
		"11000110000100111101111011010111",
		"00101111100111101010111010011001",
		"11100001100101000110010111110011",
		"11101101100001100101111111111111",
		"00101000110011001000000111100100",
		"01001111101110110100000110100011",
		"10000000101001100011110101101000",
		"10001110100111001010100000111110",
		"00011101010000110001010011100010",
		"10001110100100111100100101101101",
		"00000110110110010110110011001000",
		"10000110010111001000010110110000",
		"10001001111111111001111100110101",
		"10011011000010110001011101011011",
		"11100100101011011111110000011001",
		"01001001101000100110111111011111",
		"11001010001100111011101101010100",
		"01010011001010110101100111111000",
		"00100000000110101100010111000001",
		"11000101000011101101001011101011",
		"01000010111111010110100001001100",
		"10110000101001000011011111000001",
		"10001100110011111101011111101000",
		"11111110110010110010011011100101",
		"01010001101100111100010010110101",
		"10010110100000001001000001001110",
		"11001100100000011010010001100100",
		"00000101110101110010010111010010",
		"11010100110110001011000101011000",
		"11001000011001001011101010100100",
		"01101001110001011110101011011010",
		"11000110010001000011111000000110",
		"00010010010100010010010100101111",
		"11000101011101011000000000110010",
		"11000101011101111000111001100111",
		"01101111100011011100010001101011",
		"00110000101010111001110101011111",
		"00100000010111010010001000100000",
		"00011000101011001000110010110000",
		"10011010110101010011111100000011",
		"00001110100000001001001000010101",
		"00010100001101101011010010001000",
		"11010000010001101000100111100100",
		"01000111111010100111110101101101",
		"11000010100000110110100000110000",
		"01100010000000010100011011011111",
		"01100101000100110001000110100111",
		"00001011100010001111010110000101",
		"01000010010010111001101110000111",
		"00110011001010001010000110111111",
		"00101001110100010001010101001000",
		"01010111101110010110111111111011",
		"10011011100101101110101010110000",
		"10000111010110100010010000110101",
		"10010010010100101111111101111001",
		"10100110001000111011001101110010",
		"00111011000001000100011111110111",
		"11000110101000011011110010101111",
		"00001100101010100100001111001001",
		"00010011101111000111111010010001",
		"11100001101000000001000110100011",
		"10011100001001100010110110110000",
		"00010001001011000101001000100110",
		"11110000000000001000101000000000",
		"11111001000011001011000100001001",
		"11001001010101000000111011101100",
		"11011100000011110110110110010011",
		"00011011000110110010000000101100",
		"00001111010111010111110000011111",
		"11101111101000011110001101110000",
		"00001110101001101110011010000101",
		"00010011010100100001100111000010",
		"10001011101011111110011111010011",
		"10101000110110100011111001111111",
		"00100011110001111111110101000101",
		"10000111011111111101000011111011",
		"00110011110101001111111001001000",
		"11100000111110111001001010110011",
		"10110001100100111000101101011011",
		"10000011010110000010100101100111",
		"01010000111001101000010010101010",
		"10101100111100000111100001100101",
		"01011011101000101110010100000010",
		"10110000111010001000000110100101",
		"01101110110010101010100000111110",
		"10110011110101111010010100110000",
		"00001110011001000011101101001100",
		"11011010001111101011000011101111",
		"00110010011101100010100011101011",
		"10000101111110100000111110010001",
		"10111100101110111000111111011111",
		"01101000100000110000010000110100",
		"11000110001001001101101011010100",
		"00000110101101001111101011100011",
		"00001101011100111011110100101110",
		"11001010010101000010100100010011",
		"01100011100000011010110010101001",
		"10010100100001111011011101101010",
		"10011001101101101101000110011100",
		"11110100011101101000100110110000",
		"11011101000101110110110100100000",
		"11010001001000011001101000000000",
		"11011101000011011000000111011100",
		"00110111000110101011010101100000",
		"10001101110010101110101101010111",
		"01011010011011011011101100110010",
		"10001010000010110011101101101010",
		"11111100010110001101000011101110",
		"10000000101000011010100011110110",
		"11100000101011000111100100101100",
		"10010000011110000101111111011101",
		"01111011001100111100111011100010",
		"10010001111100010000100001010101",
		"00001011100000001001101011000010",
		"11100100101111010011100001010010",
		"00001101100101100110001011011110",
		"01100011010100011101000110010001",
		"10110111100101000011110110011010",
		"11110111111110001100110111110110",
		"00010111100001101101010010100100",
		"10101011011000010100011111011101",
		"01010011100100101101001000110101",
		"11001101101010011110111100111111",
		"01001001101000011000110011000001",
		"00000101111111001000001110111001",
		"00010000101110111110010001001111",
		"01101101000100011001011100011011",
		"10110111000011110110101010101100",
		"11100010111111111000011110101110",
		"00101100110111010011101011111100",
		"11001111000110110001110000110001",
		"00011110010011001111111101111110",
		"11100101111001111110110001001010",
		"11010011110110110001011010111001",
		"01101011110001011101100000101101",
		"01001111111001111001111001101011",
		"11100011000011111110100100101101",
		"00010000100000101010001000101000",
		"00001110100011010101111101000011",
		"10011110000101101000000011111110",
		"01001110110110100100101100110101",
		"11111001011001110001110000100000",
		"01000100010011111100101110001010",
		"10001001011010100000001101101100",
		"00010100101000000010101111000000",
		"11111110011001001111001001001101",
		"11100010110001000111100001000001",
		"00110101101111010001010011011110",
		"11011001101000001100000111100010",
		"00100011010001010111000011011100",
		"11111001010110001010100011000101",
		"11011111001001000110100011101110",
		"11101100111100101001001011101100",
		"00111101001011101100000111011111",
		"00010101000010110111011100111010",
		"00101001011111011001101101111010",
		"01010000000011001011010010001100",
		"00111111101001111011101110101101",
		"11100100010101111010001111000010",
		"11001100010011101100010101000101",
		"00011011010011111100010000011001",
		"10001010001111110100001001010100",
		"10100011110100001100010111000000",
		"11111011110110000011000110000110",
		"10101110000010110001101100111011",
		"01000100100001010011001000110001",
		"10010110111010111110101001001100",
		"01111011111001010111000000011011",
		"01111011010000101001000011010100",
		"10101000011110011110001110100101",
		"00100101111001110110010101111110",
		"10101111010000001001111101010101",
		"10111111010010110110010111000111",
		"00001111111010100000010111001111",
		"11011011001101000101000010100001",
		"01001010010000000011101110111111",
		"01001000010110111011111011111000",
		"11000011011001111101111100110001",
		"10110110000111011001101001010010",
		"00111011000110110111101100110111",
		"11001110100000101010101010101101",
		"01000101000010010010100000010001",
		"00110001000001000101010001111011",
		"01100001001110100001111101110110",
		"01110010111101110111001111000000",
		"01110010001011111101010111110100",
		"10101000011100010100110001101011",
		"10110110110010010011100011010101",
		"11010100111110011111101000000110",
		"01111111011100011000111000100110",
		"01101011111000111010110001001111",
		"00110011011110001111111000001010",
		"11001100011100010111110110110001",
		"11100010000100100110111010001001",
		"10010010010101001011111111000110",
		"00100100011111010100010101110100",
		"00001010010110011101000111000110",
		"10100000000001100111111101001110",
		"00000010000111010010000111011101",
		"11110101001100101111100100000111",
		"00111010010100111011000011111001",
		"01111010011010101101101001110000",
		"00011011000101000011111011110011",
		"11110010111001101110111001101111",
		"01000001010000011100001000011100",
		"11111000010111001001100010010101",
		"01000100110000101101001111110001",
		"00110010010100101010001011101000",
		"01101101010110001011100110111101",
		"10001100011000001010000100011101",
		"10101111111100001010011111110101",
		"01101000000010100011110111111101",
		"10010100100111010001110100001100",
		"00011101101110001101100011000101",
		"10001011110001111101101110010100",
		"11110000110111010001001110011011",
		"01011111100001110000110011110110",
		"00100101000100011001110111101001",
		"00111110111011101000000010101001",
		"11100001001110001000111011011101",
		"11001010010101000100111010000111",
		"00001110100100011011011111000011",
		"01111101101100011100010101101111",
		"10001111111000111011000100000010",
		"10001010011000000001000001110011",
		"01011101110001101111010011011110",
		"10101100100000001111100100001110",
		"00010001111100110110010101010010",
		"10000111000010011000110001101011",
		"00010100101111000100111110100110",
		"10000001111101100010001000001110",
		"11111011011001001101001111100100",
		"10111000001111000011011010010111",
		"01101100000111001100010100111010",
		"00011111001101011011111110000111",
		"01110111110011010011000010101000",
		"00011000110110100011110111000000",
		"00111111110011111000000011101100",
		"11111100000001111111011110011101",
		"11101110000000110010110000000111",
		"01100101111100011110100000001001",
		"10100000000001101001000010011101",
		"10000110101100010100111100111001",
		"00101000000010011010010100011001",
		"01000110011100101010100111110110",
		"01010101110011100010010110001000",
		"10111011101001101011010010000001",
		"11101100001000000010100011000101",
		"11010110010100000011001101110111",
		"01100000001001001111010001010100",
		"11010001011000001010110101001001",
		"01110100101101111010001101101001",
		"11111101000001011100100111111011",
		"01111010100101010110000001100110",
		"01011000110110111101001000111111",
		"11101101010110110001011110000011",
		"00001001100101101010100111101110",
		"00101111110110000010000100101000",
		"10111110000110000010101111000011",
		"01011110100111111010011110101011",
		"11011001111100001011001110111110",
		"10001001010111010001100110101001",
		"10101100010100110000010111111100",
		"01100010100111001100100001110111",
		"00001010110101000110011110010110",
		"01010010000111011011010101101110",
		"10010110000100001100111011000001",
		"11101000010010111111111110101110",
		"10110001000101101100001111001001",
		"10000110011011001101100001111001",
		"10111111001101100100011111100110",
		"11110010110110010110111000110001",
		"01110110001011010001001010111011",
		"11110011011010110100001001101001",
		"11000011001101111111011011001110",
		"01100110011110101001111000000011",
		"11101010001110111101011111101010",
		"01101001001110100010111001000000",
		"10011101010111100101111110110111",
		"00010000011110100100000101110100",
		"00101110010010000010001000000011",
		"01110011011010110000010000000010",
		"00100010001110010110111010011111",
		"11010100000010000011001100110111",
		"11000000010111011011110101000110",
		"10000010010011111100011101001101",
		"01110000111000001110110101010010",
		"10000111001100101011100110011000",
		"00101101001000111010010111111110",
		"01010011010010111110011001100110",
		"00000101001100010010110111100111",
		"11111001100101000111010100101111",
		"11001100111111101110111010001110",
		"00111000001011100000000001101110",
		"11100111001111110001101010000101",
		"01011111000001001101001101101000",
		"11010010100110100110010111100011",
		"11111100100011110110100111000010",
		"10101111011100110000000111011100",
		"11000001101110111000100100011011",
		"10010010111000010101101111010110",
		"10000011110011010011110001101001",
		"10001101010011101001110110111111",
		"00110011101010110011000101000011",
		"01100111000001010111001100100001",
		"01101101111001010001101001000101",
		"00000011110010110100101011001010",
		"00000100011111111101101110001010",
		"10101011000101100011011100001101",
		"01010100011100111110101011000101",
		"10001100111001100101101010001101",
		"00110011101011100110110101101111",
		"11000011010110000110011101111111",
		"10101011111010110101101110010010",
		"10100111001111110110110100011111",
		"00010111111010001000100110111011",
		"00111111110110111101110111011101",
		"11000100001101101010101100101101",
		"01101011001011010001001000011100",
		"01110011010010001010111001010100",
		"11000101100100101100111101001101",
		"01011000001100100111110101100011",
		"01010111001111100011011100111000",
		"00110000010000001011111011101011",
		"11101011011011101011001001000100",
		"10010010010000101101001100101011",
		"10011110000111101010000111000111",
		"10101000000001001000000011111101",
		"00010101110101100001101011000010",
		"10010011111010010011001100011101",
		"01011010100101110111101000010000",
		"10000110111001101100000000111001",
		"11110001011011010010000000011100",
		"11111100010001101101011110111110",
		"00000110000000111000010000110011",
		"00011010111100001011111001100011",
		"10101111010001001110011000001011",
		"01001001101010001110111101110110",
		"11010111000110001001011011010111",
		"01010111110110001110101000011000",
		"11101011010101011111011001010011",
		"00111101001111111110000000100100",
		"01011011011100010010111110001001",
		"11100011111100111011011100100011",
		"00100011110000110011110100011110",
		"11000100100110100011111101100110",
		"00000010010001001101010101011010",
		"11110101100001100010011111000001",
		"11000110101011110011101011111000",
		"01101011101101011000110110011100",
		"11100111000011000000111111101000",
		"11010101110001100011011100000001",
		"10110001010110000000011001110110",
		"00010111000101011000011111100000",
		"10000101100111001011111110100100",
		"00100011011000000101111001100101",
		"01101111100011001011101110100000",
		"00110111101000011101011111110110",
		"01010110000101001010011011000110",
		"11100000000010011101110110001000",
		"11100100001110100101010001010101",
		"00111111101100111011111000101000",
		"00101110111011011011011101110110",
		"11110100010111101010001011101101",
		"01100011101001000001100100111010",
		"00011111110000001101101101101111",
		"11011010101011111011010111010110",
		"11111011001100011000000010001100",
		"11110110111110011011010001010101",
		"11000000110010111010100110001100",
		"11111011100111101001100111010101",
		"01101101110100101111100010001000",
		"01010011001100101011100110011101",
		"00010000111001011111111100011111",
		"01110011010001111010110011110011",
		"00101100000110110001100101100011",
		"10111110000111100000000000001111",
		"00110111000000011110110010100111",
		"00111010010111111110001101101111",
		"00110011011011011111001011110010",
		"00110110110110100101101111000111",
		"01111011001000111101011010110110",
		"11011110011100100111100111011101",
		"01111110011110001101010110001000",
		"10110101100101100000100000011011",
		"01011111100111010111110000110010",
		"00010110001001001000010010010111",
		"00011001111010000100010010011101",
		"10000100000010111100001111000110",
		"11000010100101110011010111011001",
		"00001001001111101101001000010101",
		"11010010011011011100110000000111",
		"01000101111011110110001010110001",
		"01110111100001110011101101110011",
		"01011011001111000010100111100000",
		"00000010000000001101011000101101",
		"10110101001010011100000011000001",
		"01110111010110000011011111101101",
		"11111111000010000101010010001111",
		"10011010011000010110011001010001",
		"10001001111011001110111001000101",
		"10010100001000011110111011100100",
		"00110110100101101011011101011000",
		"11000010000000100010011000110111",
		"00011111100000100000100001010011",
		"10001100101100110100100100100000",
		"01101110011101100000110000000011",
		"11110100010000010001000011111111",
		"00001010000011100001111100111000",
		"10011000011110010100111110011111",
		"01001100111000010100000010101000",
		"11100001000111100110011001101110",
		"10001111010010101100110010000000",
		"01010101001001010101000111110100",
		"01101101011010010111001011100011",
		"00100101100101110110100001101001",
		"11101001101011011101110101111110",
		"01110011101001000110000010100011",
		"01101001011111110011100101001110",
		"11010010111011000111110110110111",
		"01010011001010011111111011010000",
		"01110000110000111111111100101010",
		"11000110001001100100000001111100",
		"00011100100100110010111011111010",
		"10000001010110100101000001000100",
		"01101100110101110000100001101100",
		"10011001001001110110110011000110",
		"11111001100010110101001101010101",
		"11100001010111011011100001001111",
		"10000110001101111110000111100110",
		"11101101010111001111101110111001",
		"10110010101101000001011100011100",
		"01101100110111100001000100111000",
		"10000100000010100011111001111010",
		"00101101001001001100101111111110",
		"10001100111110101101011110000111",
		"10100110010100001000010111011001",
		"10000000010000000011010001111000",
		"10110011111110110010110000100101",
		"10001001001011001001001110010101",
		"00111001001110000111100100101101",
		"00000101110100000110100111101010",
		"01000110011100010010000101100001",
		"01101001111001101001111101011110",
		"01001111010101110101001011111101",
		"01111011100000010100001001011010",
		"11101001111000111001011110010110",
		"01000101010111010100101101000111",
		"10110000011101111100100001000111",
		"00000101111100011100100001100111",
		"01111101100110011000111111110001",
		"00010010110011001101110110100111",
		"10001000110100001010111111000110",
		"10101000111101000011101101001110",
		"00010011101001100101101110010101",
		"01101010101011010100001101011110",
		"00001011011000010110110111000110",
		"00011001101100101000001010100100",
		"11100000001001111001110101001001",
		"11110011110111101011100010100000",
		"10001011010101011110010000101011",
		"01101101000111111010000111101111",
		"00110001100110101111001111110010",
		"10110111101110110110101000110010",
		"01100101111010101100001110110110",
		"10001001100001111010100001101010",
		"10000011011011110010000011000011",
		"11011110000101111010011110111010",
		"00011010001101101001011010010110",
		"11111110101011101000110011101111",
		"10011101110000111000100111110000",
		"11001001000110001001100000101001",
		"00000101000001000010110111100110",
		"11000001101001100001011011101110",
		"01111011001010100101110110010100",
		"01001010000110001011000011000011",
		"10000010111100110110000110010011",
		"11101101110011001011111001111001",
		"00001000101101100001010110010110",
		"00010000110100011010010001000010",
		"00001100000100101011011101001010",
		"10001010110010101001100001010110",
		"11010101000001100001001111010110",
		"00011010110010001100110011010111",
		"11011001101111011110100001111011",
		"11011101100110000100001100010011",
		"00101111111101100001000001100101",
		"10101101100110010110111101001011",
		"10100110010000110111000100100011",
		"11110110001100100111101101000001",
		"10011011011111001000000000111001",
		"10010101111110001010000000011011",
		"00111111000011011010111110011111",
		"11011110110001100001111110101110",
		"01010111100011010010111110111000",
		"10111100111000101000011100011101",
		"01111110111000100011100000000100",
		"11000110001111101011100110010010",
		"01000011001111011101100000111100",
		"10000010011101110111001101001110",
		"01111110000101001001010001101010",
		"10111100001100011010101111011001",
		"01001111001111010110110100101110",
		"11101110000011101100111000111010",
		"11010000010001001100010011000010",
		"11111110101000000111101100110111",
		"11010010110000000010101010001111",
		"10001101011000111101101001000111",
		"00010001111101100011011001000110",
		"00001001110010110000111111001001",
		"10110110101010000101010011101100",
		"11001100111110000100000011010110",
		"11000100110110100111111101011100",
		"10110010110011101100110110010110",
		"11111101111101110011110000100111",
		"01101101010110011000111010100101",
		"01101001011110100001010101110011",
		"01110111100101111000100001011110",
		"01101110101110110010100000000101",
		"01000111110000101110100111001011",
		"11111011001001011111110110011101",
		"00000100100001101011111100101111",
		"10001101010011011100111011110000",
		"00010101100011101110110011010110",
		"10011111100000100011110110101111",
		"01100101111100110011110110110010",
		"11110111111001010001001010101100",
		"00101001100010000010001000101101",
		"11000111100101010111011111101110",
		"01100001011110101110111110101100",
		"10010100111100011101100100000110",
		"11101011000110101100011001100100",
		"00101011100101010001000100000000",
		"01101110000110110111101001000110",
		"10111000010010010011011111101101",
		"11000010111010101010110011100110",
		"01000010010011010000110111101110",
		"00000000001010110000101110000000",
		"11011011111101100000110100011001",
		"00011100100011110010010101001101",
		"00011000010001101110100101101010",
		"01001110011000101101111011111101",
		"10001011100000100110110111001001",
		"01101000000110111010000100110011",
		"01111110011110000001001100101101",
		"00100001111001100010111010100110",
		"01110001100101011101001001111011",
		"11110101100011101100000110111010",
		"10101110000001111010111010111111",
		"01011001101010111000111101110011",
		"10100000001100101110101010111010",
		"01111010101000000111011000111100",
		"10100100011110010100011011001011",
		"10110111100000101001100111011100",
		"10110101101100100010110101100110",
		"11010111110111101101001100001011",
		"10110010100111000101101010010000",
		"11111000110010001110010110011101",
		"11010001011010011111111101000110",
		"10100110100101001110101001000001",
		"00001001110000011001001111010011",
		"00001000000001010110101000111000",
		"11000011001111101110000001111011",
		"11001101101011000010001111101100",
		"01001100100011001010010110010110",
		"00001010010110010101100101001110",
		"10110011010111111011110000101000",
		"10111011111100101001001100100001",
		"10011010001101101001011101100101",
		"00000110000010100110100001100010",
		"10010011011010011010100100100000",
		"10101000100111101001011101011100",
		"10100110000001101111100010110000",
		"11100101111100101010000000010000",
		"11101011010010011000100100001100",
		"01000110111011100110000100001110",
		"01011101010011100000000010001111",
		"01000111111110011001100001001100",
		"01110000010101101001011001111001",
		"10111001010001010010001001011110",
		"00000000101001011001001000011100",
		"10110001000101100011111101000111",
		"01110001100101111111111100101011",
		"01111110011101000010010011110010",
		"11111111010011010000000111001000",
		"11001100100111110111111110000010",
		"10010100011111111100011011011110",
		"11000110100110010101111111000000",
		"11101001001110100111010101100101",
		"10001010101110000000011110100111",
		"01101010100110111000000111111100",
		"00001101110010101100001100010001",
		"01110110111111100001011010111110",
		"00011111111111000001111100111100",
		"00110101001111101001010100111000",
		"10111100100011001110001101011010",
		"10001001000011110111011010110010",
		"11111110010100110010011001001110",
		"11111100111111110101111010001001",
		"11101100001111101101010111110000",
		"00001101110001001001101111100101",
		"01101010011011010101100001001101",
		"11001000110101110000011111101110",
		"01110110101110101110000101101001",
		"10111111001111110011111001011010",
		"01001011001000100000011001101110",
		"11001010010111000111011001010111",
		"10100001000100011111111110011101",
		"11111101011111100101000100011001",
		"01110000011011110110100101011110",
		"11111000001011111011100011110111",
		"01011000110101110101111111111010",
		"10010011111001010111100111001001",
		"10001010110001101101010110011001",
		"00010110101011010001101011000100",
		"01000111100100111111011101101111",
		"01111000100101000000001001111000",
		"00001000101010001010111111101010",
		"01110000101010111110110111011110",
		"11000000000100101010111010001001",
		"00001001110101110001100101111110",
		"11011011111001001111000000000010",
		"01011111110100001010000110010101",
		"00110111100101001011010110001011",
		"10010010010101010001000111010001",
		"10101011111010010010100111011010",
		"11011000011101001100111110000011",
		"11001000100111111000110001010110",
		"10001110111001000000100011110001",
		"01011000101101000111011110111000",
		"10001111011110110111010101100110",
		"10010001000111000000100000000100",
		"10010010100110010111101010100100",
		"01101100110110100010001101100011",
		"11111010101111100010111101100101",
		"00010100011001100010110101100001",
		"00010110101011001001001101010010",
		"11010011001000011111110111101100",
		"10110100000001111011001101110010",
		"00000110111001101100110100111101",
		"01000110101000010000010000101111",
		"00001000001001110000111110010010",
		"11111000000000011010011010001101",
		"11111001011110011110001001011010",
		"11001011001000110000001010111010",
		"00101011011011100001011010101001",
		"01001000000110101111010100011111",
		"11111011101011001010001000110010",
		"01001001001011001100111111000110",
		"10111110001101110101111100011000",
		"00101000011100001010001000100110",
		"01111000001110001100100011011000",
		"10001011011011110000101000111110",
		"00101101001111111110101101000111",
		"00000100000001011011001110001101",
		"11010010001000011111101101110000",
		"10110001100111010010110100101110",
		"01000110010011001010001111101000",
		"10000001100010100010001101010110",
		"00010101101101010110010110000111",
		"11110111010001001011001001111110",
		"01001010010010111010011101000101",
		"11000000000000011001011000000101",
		"00011100110100010110001110101010",
		"00101110010111110001110000111111",
		"11101111110000001000101100100011",
		"00110001010000101001111101011110",
		"10100010111110110000001110001110",
		"10010100000011101111000010110001",
		"11101100111110010111101110001001",
		"11001010011101110001111110001111",
		"01010000001000010010110110101011",
		"11110100101010101110000000110010",
		"01010001110110101100010111110000",
		"11011001110011010010011101000100",
		"01110001001100111110000010100010",
		"10101101010100110110110101111010",
		"11001101001000101110010110110011",
		"10100111110100100010101101010100",
		"01000111000001001101001010100001",
		"01101000111000110011101001010100",
		"00011011011110110011011001100011",
		"01010101001011100101001100100011",
		"10111100001100101100100101010110",
		"00100011110011001101101110011111",
		"00010111100010001010110011101101",
		"00011011111110100101111100110101",
		"00101111001010000111101101111111",
		"11000111101001001010001011111111",
		"01011110010001000010101001001011",
		"11101010001011011101011000000000",
		"01110000000100111111111010011010",
		"10001001101100011111100101011000",
		"10111111111001100110100110010010",
		"01101000111101110100011011011010",
		"11100011111101001100101100001101",
		"11110111001110101011110001100101",
		"00111100010100000011100000110011",
		"10001100001101101111001100111000",
		"11010010011100110000111000011100",
		"01000001111101101101101110111010",
		"01111100000011100000001011100000",
		"10100111011001111110101111011111",
		"01100010011000011100001100010000",
		"00101101000010111001000010000111",
		"01110100101001010001010000000010",
		"01110010101110011110001010100101",
		"01000001100011010111100000111001",
		"10010010010110100101100111010101",
		"01001101100000111011110001100101",
		"00111110111001011101011011101010",
		"00100000001001011111101110100110",
		"11001001000101101101101111101100",
		"11110110001010001101111110111110",
		"11111111110011100000011011100111",
		"11011100001100101000101101100111",
		"00010101100110000100011111111000",
		"00001010010010100111101100110110",
		"11001000101000100101001110000001",
		"01100011100010100011101100100010",
		"00101001111010101101110010100010",
		"01011100001100101100011001100111",
		"00100100101010110100000111001001",
		"10100110100000010011011100100000",
		"10000011001110010101001011011001",
		"10110101000001001101000110010111",
		"10110000101001101110101000111111",
		"10001101000110000000010100010011",
		"10111011000110101100010110111011",
		"00011110001111000111010010100010",
		"00110111101001110111111111011000",
		"10110000011100010100001100011100",
		"00101000100010010110101111101100",
		"10110011100110100000010000101110",
		"10110000100100110111000000110000",
		"00000110000101001111110100001110",
		"00001110011111010101001000000100",
		"10011000000100011100010101101100",
		"01110010010100110100101001000001",
		"00011100010100010101011111100110",
		"11100101101010010001011110001100",
		"11010101110111101011010101100001",
		"11000100111010010111110100001010",
		"00110110001101110000111000001101",
		"01111010000110011000011111000111",
		"10001010010100010100010101101110",
		"10110010011001100111100010111011",
		"01000010111000101001011011001000",
		"10000110000110000001010101101010",
		"01011111111011111011001000111111",
		"00011100000101010100000010100000",
		"01000101001100101000011101010100",
		"01111010110100010011011001111110",
		"10110000111011010110110001100010",
		"00011010010011101000111100110010",
		"11010000001100111011011101110101",
		"10111010011110001100111101000010",
		"11111110110110110011011001100001",
		"11110100010100010101000010010111",
		"01111011111100001011011011111111",
		"01111011001010110010000101110101",
		"11110100011010101010011011111001",
		"10100000100011110100000110101001",
		"11111011011100101000010101000110",
		"10100001010111010000011001110000",
		"11010111100100101111000001100010",
		"10010001110011000000100010001111",
		"00110110111011000100100011111100",
		"10101100101001011110010010101010",
		"11111110000011011000011101001101",
		"11100010110100000001110000110100",
		"10011111011011111100011101000110",
		"11100010110111001011100111100111",
		"01010000101110100000001011001111",
		"11000100011000000010111001000010",
		"11001000000011000011101110101100",
		"00111110101110010101111011000011",
		"01000000001110001011010111111111",
		"10010001011111010101111001100110",
		"11000011000011110111001011101111",
		"10010001000000000110010110111110",
		"11001110111010111101110001110110",
		"00110011010100000000111001110011",
		"01111111110011000110000111111001",
		"01011100111010100001101010110011",
		"01110010110111111110111111101111",
		"01011110111110010000010010001011",
		"10110000111100001010100001001001",
		"10101000100011100000010000000110",
		"00101010110101011010111101010010",
		"10101010011100000110100001100011",
		"00110101011100100011110101001101",
		"00111001010010101111101000010100",
		"10101011110111110111100011010101",
		"01011001001100001011100110100001",
		"00111010001000100100001010010111",
		"00001100111100110010100111001100",
		"11100101111010110011100010000100",
		"10111011101111011001101101000101",
		"00010010000000101000010110010010",
		"01110110000001101111000101001010",
		"10110100010111000011000011110001",
		"01001110100100001101111110100001",
		"11110111111011110000101001011101",
		"11011001001111011101011100101110",
		"10101011000001011101011100000110",
		"01011000111100100101101111111000",
		"11010101101001111000101000101000",
		"10011100011100111001010111101010",
		"01110000100010110001001000010001",
		"01101101000000011100010101011110",
		"10110100101111011001100101101110",
		"11011000010100010101001001001101",
		"00111111011110110110011011100101",
		"00111100111010100011100101101100",
		"10111100100010010011001111010101",
		"01001011000101010100001110111101",
		"00011011010000010001001011101010",
		"01110010100000111011011011111101",
		"11011110100001011111011101110011",
		"01101000101111101000010011111001",
		"01000111000111001000111010010100",
		"10010011111111101010110010010001",
		"11010001100000001111100101110001",
		"01110010110001010100110110001011",
		"11111101001010100100011101111000",
		"01010111111100001010011010111111",
		"01110101110001101100000000011000",
		"10000011001001001110101001010000",
		"00110000001100000011000100010011",
		"11000010110101100100101111111011",
		"00011110110000111001111000000110",
		"00010111010010111110010001000111",
		"00111100001111011100000101011110",
		"01111111010100110101100100000010",
		"10001001101001000001100011010101",
		"01110000010100100011100011100000",
		"11000010111001001110000010101000",
		"00011001011010100001010011110001",
		"00100000010010000110000010101101",
		"10001101011010110110110010111101",
		"11111100001110101100100110000011",
		"10110111001101111011110011111000",
		"10010010101001100110001111101000",
		"01000001110011010001110101100011",
		"01100101001001110100101011000100",
		"01101111111000010011111111001010",
		"11100110001010101000011000010110",
		"00110010110011011011011110101001",
		"01111101011110100111100000010011",
		"10101000001011100001100101101100",
		"10001101100101001100110110001010",
		"01001100011001110101001101010100",
		"01010011000010011100101000011111",
		"01110010110001010110011010011000",
		"00100100100110010000111111010011",
		"00110001011110110010010011011110",
		"10001000101011011110101101110100",
		"01011100011001110010110001111100",
		"01111010111000111100101101100110",
		"11110110111101101011100101111110",
		"00100110110110111001110000011101",
		"10010000100010011001110101011011",
		"00110101100100010010111001110110",
		"10111011010100011010001001110000",
		"01011011110000101000111111011010",
		"10000100000100000101101001100001",
		"01101000000000110110111111011011",
		"01101101111100001011100110011101",
		"00001101100111001010101100100010",
		"10010010001010000110011111101001",
		"11010100011000100100011100011010",
		"01011111000110000010111001001001",
		"01101010001010000011001010001110",
		"11100110111000100010011101110111",
		"01111111100000001001011010111000",
		"01100011001110111100110011001010",
		"01100001010100101000111000000101",
		"11001010000110011110111110110000",
		"10110010000011000101100100000010",
		"01111000010100111001100101010110",
		"10111001101101010111001100011001",
		"01110101111000001100010011000001",
		"10110111101011110111011011001100",
		"11000000011111101001010101010110",
		"01101100110011111000011110101111",
		"10010110011111000100100111000011",
		"01000000000011010100100001011000",
		"01000000001101110011111011011000",
		"00111001101000100101011010101101",
		"11001000001010010010111001000101",
		"00100011111001100010000111111000",
		"10001111011010111010110101110110",
		"10110000000111011010100100000110",
		"11100110000101111100100010010011",
		"11101010001010000111011010111010",
		"10100110111110100111100100000001",
		"00110101100000110100100010001001",
		"11100001010010001010000100011111",
		"10111101111111011111101000010110",
		"01011101010111100000101100110001",
		"10101010011101000101001010100001",
		"01000101000101110000111011011010",
		"00100010000000001100110100001110",
		"00000011001011100001000011111001",
		"01010001111010111011100010000100",
		"11011101011001001110001001110011",
		"11011110110010111100111010111000",
		"10000111001000000100110001100111",
		"00000001101111000011001110011001",
		"11110110010101001111110101010001",
		"00110110101110110100111101000111",
		"01110100010001001111000010111111",
		"11010000001100010111000010010001",
		"01011111110111001010101011000011",
		"01011100110011011010000001011011",
		"00011111000100101100111110000001",
		"00111111111011111100111010111010",
		"11001100011101010001111010010110",
		"11001001101101010110010100011001",
		"10111010011011011101011110000101",
		"11000110010000101100111010100000",
		"10100111000101110100111010010001",
		"01010100111001100100010110100000",
		"00101001100000100000111100111101",
		"00010111111111000101010001001000",
		"00100100000111110011101000111010",
		"10100000110101000101011110101110",
		"10111101011111001100000110001000",
		"00000001011001110100000100101110",
		"00010111110110100011101010001000",
		"01110001001001011110001110000000",
		"11111010010101001110101100011110",
		"00001110110000000011101011111100",
		"01001001110011101000010101100011",
		"00101001111101001000101000011010",
		"10100001100101011010001101101011",
		"00010100100011111100101101000001",
		"00000100100010111110011100111000",
		"00011100000011100100011001010001",
		"10000110010010100100101000111111",
		"01100010000110000100010110001010",
		"11011001111101100001011100000110",
		"01110001111101001000111001101100",
		"01000010010110001111100110111100",
		"11010011111011010111010001100011",
		"11000010100000001001010110001111",
		"01000000000010101110010001101010",
		"10011000111111101001101001000101",
		"10001110111011010101000011111001",
		"11001010101000011011011111111000",
		"01110100000101110100111101111000",
		"00111000100011001001001001011010",
		"11100011000001101001011111110011",
		"10011110001100100010001110101110",
		"10001101010000110100010000100111",
		"10001101000100111100111010111001",
		"00010110010101010100000000001111",
		"00000010111000100011101100000101",
		"10010010001100100110011111100110",
		"01101101000010100000001100101011",
		"10011100111101101100011111111010",
		"10000110100001100010000001001100",
		"11100111100011110111000010010101",
		"00001101111011101001110010010001"
	);
	signal clk                : std_logic := '0';
	signal rng_ce             : std_logic := '0';
	signal rng_mode           : std_logic := '0';
	signal rng_s_in           : std_logic := '0';
	signal rng_s_out          : std_logic := '0';
	signal rng_r              : OutputType;
	signal rng_s_out_buff     : std_logic; -- need to buffer in a register ourselves
	signal readback           : StateType;
	constant initState        : StateType := "1010100010011101101011010011101111100010001111111100100101011001001100110000001111000101011010111100010110011000011110001101000010010111110010010011001001111110010111100110100010100101000110010101111111101111110011001000011010101111101001101000001010111010110111111101000010010010001001001110100100111011001010000111111111011111111001110001001100011111010010000010010110111110100010111011111001010111000110010010000000001011000011011001011101001110010000110001011110110001110010011000110000110000010100001110110110000000000110111101010000101111000000100101100011011111011100011110000001011110000001001000100010101011010010010101100101111001001100011010011100111110101111100101011000111100010011110001110011110100100011110010111101100000100010011010010111100011010110000100011000101011111110010111110111110100100110011101101010101011001000100110100101010000100100110011011010100110010110010011100100111111010110101100010000111011001011001011100100111111110100001000101011000111110001100000100111001100011010010111110000010110";
	constant refReadback      : StateType := "0100000111000111000100000011100001101010010110011001010010000000101111000100011101100101100101111010001010110100100100011110000110011100100000001001110110011111001001001001101000001100111101000011111111001000001011101101100011111101001100011101011100000100100011110111010011110011101100001110011010111101101101101011011100000101000010010001100100101011000101010010110010010110010100001010010000001011001111111000000101000111010111100001110011100011101111111101111010011000010111110000100001101110111010000000010010101011100010101011001111100001100101111010001101100001101101000100100000011100000001010000110011111100111100101000000001111000101001000010011010111011000011111011101000010011111000010001110010011001110011001100111001100000011001101000001111111010100010110110110010001101000000010110000011100000111001111011101011100101011001010011010110011101110110001000110011000100010010110000010100001111010111110100001101111110110110011101100000101011101000000100101100010001110010110000001000111100011011000101011001110101";
begin
	-- Instantiate random-number generator
	uut: entity makestuff.rng
		port map (
			clk              => clk,
			ce               => rng_ce,
			mode             => rng_mode,
			s_in             => rng_s_in,
			s_out            => rng_s_out,
			rng              => rng_r
		);

	-- Drive clock
	clk <= not clk after 5 ns;
  
	s_out_buff: process
	begin
		wait until rising_edge(clk);
		rng_s_out_buff <= rng_s_out;
	end process;

	tb_driver: process
	begin
		--First cycle of state loading
		wait until rising_edge(clk);
		rng_ce <= '1';
		rng_mode <= '1';
		rng_s_in <= initState(0);
		
		-- Continue loading state
		for i in 1 to N-1 loop
			wait until rising_edge(clk);
			rng_s_in <= initState(i);
		end loop;
		
		-- Switch to rng mode
		wait until rising_edge(clk);
		rng_mode <= '0';
		
		-- Here the checker is looking at the output
		for i in 1 to 2*N-1 loop
			wait until rising_edge(clk);
		end loop;
       
		-- Start reading (and loading) state
		wait until rising_edge(clk);
		rng_mode <= '1';
		rng_s_in <= '1';

		-- Continue reading state
		for i in 1 to N-1 loop
			wait until rising_edge(clk);
		end loop;
	end process;

	tb_checker: process
	begin
		wait until rising_edge(clk);
		wait until rising_edge(clk);

		-- Wait while state is loaded
		for i in 0 to N-1 loop
			wait until rising_edge(clk);
		end loop;

		-- Check output over following 2*N cycles
		for i in 0 to 2*N-1 loop
			wait until rising_edge(clk);
			assert rng_r = expectedArray(i) report "Output mismatch." severity failure;
		end loop;

		-- Read state over N cycles
		for i in 0 to N-1 loop
			wait until rising_edge(clk);
			readback(i) <= rng_s_out_buff;
		end loop;

		wait until rising_edge(clk);
		assert readback = refReadback report "Readback state mismatch" severity failure;

		std.env.stop(0);
	end process;
end architecture;
