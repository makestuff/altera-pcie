--
-- Copyright (C) 2014, 2017 Chris McClelland
--
-- Permission is hereby granted, free of charge, to any person obtaining a copy of this software
-- and associated documentation files (the "Software"), to deal in the Software without
-- restriction, including without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to permit persons to whom the
-- Software is furnished to do so, subject to the following conditions:
--
-- The above copyright  notice and this permission notice  shall be included in all copies or
-- substantial portions of the Software.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR IMPLIED, INCLUDING
-- BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND
-- NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM,
-- DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
-- OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE SOFTWARE.
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library makestuff;
use makestuff.util_pkg.all;

entity util_pkg_tb is
end entity;

architecture behavioural of util_pkg_tb is
begin
	process
		procedure test_log2(
			constant value    : in natural;
			constant expected : in natural
		) is
			constant result   : natural := log2(value);
		begin
			assert result = expected report
				"Expected " & natural'image(expected) & " from log2(" & natural'image(value) &
				") but got " & natural'image(result) & "!"
				severity failure;
		end procedure;
	begin
		-- Test plan generated by this bit of Python (with a fix: log2(536870912) should be 29, not 30):
		-- #!/usr/bin/python
		-- import math
		-- for i in range(2, 35):
		--   print("\t\ttest_log2(%d, %d);" % (i, int(math.ceil(math.log(i, 2)))));
		-- for j in range(6, 31):
		--   for i in range(-1, +3):
		--     val = int(math.pow(2, j) + i)
		--     print("\t\ttest_log2(%d, %d);" % (val, int(math.ceil(math.log(val, 2)))));
		--
		test_log2(1, 1);  -- wrong, but more useful than making log2(1) == 0
		test_log2(2, 1);
		test_log2(3, 2);
		test_log2(4, 2);
		test_log2(5, 3);
		test_log2(6, 3);
		test_log2(7, 3);
		test_log2(8, 3);
		test_log2(9, 4);
		test_log2(10, 4);
		test_log2(11, 4);
		test_log2(12, 4);
		test_log2(13, 4);
		test_log2(14, 4);
		test_log2(15, 4);
		test_log2(16, 4);
		test_log2(17, 5);
		test_log2(18, 5);
		test_log2(19, 5);
		test_log2(20, 5);
		test_log2(21, 5);
		test_log2(22, 5);
		test_log2(23, 5);
		test_log2(24, 5);
		test_log2(25, 5);
		test_log2(26, 5);
		test_log2(27, 5);
		test_log2(28, 5);
		test_log2(29, 5);
		test_log2(30, 5);
		test_log2(31, 5);
		test_log2(32, 5);
		test_log2(33, 6);
		test_log2(34, 6);
		test_log2(63, 6);
		test_log2(64, 6);
		test_log2(65, 7);
		test_log2(66, 7);
		test_log2(127, 7);
		test_log2(128, 7);
		test_log2(129, 8);
		test_log2(130, 8);
		test_log2(255, 8);
		test_log2(256, 8);
		test_log2(257, 9);
		test_log2(258, 9);
		test_log2(511, 9);
		test_log2(512, 9);
		test_log2(513, 10);
		test_log2(514, 10);
		test_log2(1023, 10);
		test_log2(1024, 10);
		test_log2(1025, 11);
		test_log2(1026, 11);
		test_log2(2047, 11);
		test_log2(2048, 11);
		test_log2(2049, 12);
		test_log2(2050, 12);
		test_log2(4095, 12);
		test_log2(4096, 12);
		test_log2(4097, 13);
		test_log2(4098, 13);
		test_log2(8191, 13);
		test_log2(8192, 13);
		test_log2(8193, 14);
		test_log2(8194, 14);
		test_log2(16383, 14);
		test_log2(16384, 14);
		test_log2(16385, 15);
		test_log2(16386, 15);
		test_log2(32767, 15);
		test_log2(32768, 15);
		test_log2(32769, 16);
		test_log2(32770, 16);
		test_log2(65535, 16);
		test_log2(65536, 16);
		test_log2(65537, 17);
		test_log2(65538, 17);
		test_log2(131071, 17);
		test_log2(131072, 17);
		test_log2(131073, 18);
		test_log2(131074, 18);
		test_log2(262143, 18);
		test_log2(262144, 18);
		test_log2(262145, 19);
		test_log2(262146, 19);
		test_log2(524287, 19);
		test_log2(524288, 19);
		test_log2(524289, 20);
		test_log2(524290, 20);
		test_log2(1048575, 20);
		test_log2(1048576, 20);
		test_log2(1048577, 21);
		test_log2(1048578, 21);
		test_log2(2097151, 21);
		test_log2(2097152, 21);
		test_log2(2097153, 22);
		test_log2(2097154, 22);
		test_log2(4194303, 22);
		test_log2(4194304, 22);
		test_log2(4194305, 23);
		test_log2(4194306, 23);
		test_log2(8388607, 23);
		test_log2(8388608, 23);
		test_log2(8388609, 24);
		test_log2(8388610, 24);
		test_log2(16777215, 24);
		test_log2(16777216, 24);
		test_log2(16777217, 25);
		test_log2(16777218, 25);
		test_log2(33554431, 25);
		test_log2(33554432, 25);
		test_log2(33554433, 26);
		test_log2(33554434, 26);
		test_log2(67108863, 26);
		test_log2(67108864, 26);
		test_log2(67108865, 27);
		test_log2(67108866, 27);
		test_log2(134217727, 27);
		test_log2(134217728, 27);
		test_log2(134217729, 28);
		test_log2(134217730, 28);
		test_log2(268435455, 28);
		test_log2(268435456, 28);
		test_log2(268435457, 29);
		test_log2(268435458, 29);
		test_log2(536870911, 29);
		test_log2(536870912, 29);  -- manual fix 30->29 due to Python FP error
		test_log2(536870913, 30);
		test_log2(536870914, 30);
		test_log2(1073741823, 30);
		test_log2(1073741824, 30);
		test_log2(1073741825, 31);
		test_log2(1073741826, 31);
		test_log2(2147483647, 31);
		wait for 10 ns;
		std.env.stop(0);
	end process;
end architecture;
